VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO stc0_core
  CLASS BLOCK ;
  FOREIGN stc0_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1088.735 BY 1099.455 ;
  PIN ARstb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END ARstb
  PIN ClkIngress
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END ClkIngress
  PIN ED[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1084.735 916.000 1088.735 916.600 ;
    END
  END ED[0]
  PIN ED[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1084.735 549.480 1088.735 550.080 ;
    END
  END ED[1]
  PIN ED[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1084.735 182.960 1088.735 183.560 ;
    END
  END ED[2]
  PIN ED[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.370 1095.455 1020.650 1099.455 ;
    END
  END ED[3]
  PIN ED[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 1095.455 748.330 1099.455 ;
    END
  END ED[4]
  PIN ED[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 1095.455 612.170 1099.455 ;
    END
  END ED[5]
  PIN ED[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 1095.455 476.010 1099.455 ;
    END
  END ED[6]
  PIN ED[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 1095.455 339.850 1099.455 ;
    END
  END ED[7]
  PIN EValid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.210 1095.455 884.490 1099.455 ;
    END
  END EValid
  PIN ID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 1095.455 203.690 1099.455 ;
    END
  END ID[0]
  PIN ID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 1095.455 67.990 1099.455 ;
    END
  END ID[1]
  PIN ID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1037.720 4.000 1038.320 ;
    END
  END ID[2]
  PIN ID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 915.320 4.000 915.920 ;
    END
  END ID[3]
  PIN ID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.200 4.000 671.800 ;
    END
  END ID[4]
  PIN ID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.800 4.000 549.400 ;
    END
  END ID[5]
  PIN ID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END ID[6]
  PIN ID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END ID[7]
  PIN IValid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 793.600 4.000 794.200 ;
    END
  END IValid
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1088.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1088.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1088.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1088.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1088.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1088.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1088.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1088.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1088.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1088.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1088.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1088.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1088.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1088.240 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 945.940 10.880 947.540 1088.000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 792.340 10.880 793.940 1088.000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.740 10.880 640.340 1088.000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 1088.000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 1088.000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 1088.000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 1088.000 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1022.740 10.880 1024.340 1088.000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 869.140 10.880 870.740 1088.000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 715.540 10.880 717.140 1088.000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.940 10.880 563.540 1088.000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 1088.000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 1088.000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 1088.000 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 949.240 10.880 950.840 1088.000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 795.640 10.880 797.240 1088.000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 642.040 10.880 643.640 1088.000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 488.440 10.880 490.040 1088.000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 1088.000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 1088.000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 1088.000 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1026.040 10.880 1027.640 1088.000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 872.440 10.880 874.040 1088.000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 718.840 10.880 720.440 1088.000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 565.240 10.880 566.840 1088.000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.640 10.880 413.240 1088.000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 1088.000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 1088.000 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 952.540 10.880 954.140 1088.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 798.940 10.880 800.540 1088.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 645.340 10.880 646.940 1088.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 491.740 10.880 493.340 1088.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 1088.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 1088.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 1088.000 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1029.340 10.880 1030.940 1088.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 875.740 10.880 877.340 1088.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 722.140 10.880 723.740 1088.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 568.540 10.880 570.140 1088.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 414.940 10.880 416.540 1088.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 1088.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 1088.000 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1083.615 1088.085 ;
      LAYER met1 ;
        RECT 5.520 10.640 1083.675 1088.240 ;
      LAYER met2 ;
        RECT 6.530 1095.175 67.430 1095.455 ;
        RECT 68.270 1095.175 203.130 1095.455 ;
        RECT 203.970 1095.175 339.290 1095.455 ;
        RECT 340.130 1095.175 475.450 1095.455 ;
        RECT 476.290 1095.175 611.610 1095.455 ;
        RECT 612.450 1095.175 747.770 1095.455 ;
        RECT 748.610 1095.175 883.930 1095.455 ;
        RECT 884.770 1095.175 1020.090 1095.455 ;
        RECT 1020.930 1095.175 1081.360 1095.455 ;
        RECT 6.530 10.640 1081.360 1095.175 ;
      LAYER met3 ;
        RECT 4.000 1038.720 1084.735 1088.165 ;
        RECT 4.400 1037.320 1084.735 1038.720 ;
        RECT 4.000 917.000 1084.735 1037.320 ;
        RECT 4.000 916.320 1084.335 917.000 ;
        RECT 4.400 915.600 1084.335 916.320 ;
        RECT 4.400 914.920 1084.735 915.600 ;
        RECT 4.000 794.600 1084.735 914.920 ;
        RECT 4.400 793.200 1084.735 794.600 ;
        RECT 4.000 672.200 1084.735 793.200 ;
        RECT 4.400 670.800 1084.735 672.200 ;
        RECT 4.000 550.480 1084.735 670.800 ;
        RECT 4.000 549.800 1084.335 550.480 ;
        RECT 4.400 549.080 1084.335 549.800 ;
        RECT 4.400 548.400 1084.735 549.080 ;
        RECT 4.000 428.080 1084.735 548.400 ;
        RECT 4.400 426.680 1084.735 428.080 ;
        RECT 4.000 305.680 1084.735 426.680 ;
        RECT 4.400 304.280 1084.735 305.680 ;
        RECT 4.000 183.960 1084.735 304.280 ;
        RECT 4.000 183.280 1084.335 183.960 ;
        RECT 4.400 182.560 1084.335 183.280 ;
        RECT 4.400 181.880 1084.735 182.560 ;
        RECT 4.000 61.560 1084.735 181.880 ;
        RECT 4.400 60.160 1084.735 61.560 ;
        RECT 4.000 10.715 1084.735 60.160 ;
      LAYER met4 ;
        RECT 165.895 61.375 174.240 1051.105 ;
        RECT 176.640 61.375 177.540 1051.105 ;
        RECT 179.940 61.375 180.840 1051.105 ;
        RECT 183.240 61.375 184.140 1051.105 ;
        RECT 186.540 61.375 251.040 1051.105 ;
        RECT 253.440 61.375 254.340 1051.105 ;
        RECT 256.740 61.375 257.640 1051.105 ;
        RECT 260.040 61.375 260.940 1051.105 ;
        RECT 263.340 61.375 327.840 1051.105 ;
        RECT 330.240 61.375 331.140 1051.105 ;
        RECT 333.540 61.375 334.440 1051.105 ;
        RECT 336.840 61.375 337.740 1051.105 ;
        RECT 340.140 61.375 404.640 1051.105 ;
        RECT 407.040 61.375 407.940 1051.105 ;
        RECT 410.340 61.375 411.240 1051.105 ;
        RECT 413.640 61.375 414.540 1051.105 ;
        RECT 416.940 61.375 481.440 1051.105 ;
        RECT 483.840 61.375 484.740 1051.105 ;
        RECT 487.140 61.375 488.040 1051.105 ;
        RECT 490.440 61.375 491.340 1051.105 ;
        RECT 493.740 61.375 558.240 1051.105 ;
        RECT 560.640 61.375 561.540 1051.105 ;
        RECT 563.940 61.375 564.840 1051.105 ;
        RECT 567.240 61.375 568.140 1051.105 ;
        RECT 570.540 61.375 635.040 1051.105 ;
        RECT 637.440 61.375 638.340 1051.105 ;
        RECT 640.740 61.375 641.640 1051.105 ;
        RECT 644.040 61.375 644.940 1051.105 ;
        RECT 647.340 61.375 711.840 1051.105 ;
        RECT 714.240 61.375 715.140 1051.105 ;
        RECT 717.540 61.375 718.440 1051.105 ;
        RECT 720.840 61.375 721.740 1051.105 ;
        RECT 724.140 61.375 788.640 1051.105 ;
        RECT 791.040 61.375 791.940 1051.105 ;
        RECT 794.340 61.375 795.240 1051.105 ;
        RECT 797.640 61.375 798.540 1051.105 ;
        RECT 800.940 61.375 865.440 1051.105 ;
        RECT 867.840 61.375 868.740 1051.105 ;
        RECT 871.140 61.375 872.040 1051.105 ;
        RECT 874.440 61.375 875.340 1051.105 ;
        RECT 877.740 61.375 942.240 1051.105 ;
        RECT 944.640 61.375 945.465 1051.105 ;
  END
END stc0_core
END LIBRARY

