VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO lfsr32
  CLASS BLOCK ;
  FOREIGN lfsr32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN ARstb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 196.000 100.190 200.000 ;
    END
  END ARstb
  PIN Clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END Clk
  PIN LFSR0out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END LFSR0out
  PIN LFSR1in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END LFSR1in
  PIN LFSR1out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END LFSR1out
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END io_oeb[4]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 187.680 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 187.680 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 187.680 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 187.680 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 187.680 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 187.680 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 187.680 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 187.680 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 187.680 ;
    END
  END vssa2
  OBS
      LAYER nwell ;
        RECT 5.330 183.545 194.310 186.375 ;
        RECT 5.330 178.105 194.310 180.935 ;
        RECT 5.330 172.665 194.310 175.495 ;
        RECT 5.330 167.225 194.310 170.055 ;
        RECT 5.330 161.785 194.310 164.615 ;
        RECT 5.330 156.345 194.310 159.175 ;
        RECT 5.330 150.905 194.310 153.735 ;
        RECT 5.330 145.465 194.310 148.295 ;
        RECT 5.330 140.025 194.310 142.855 ;
        RECT 5.330 134.585 194.310 137.415 ;
        RECT 5.330 129.145 194.310 131.975 ;
        RECT 5.330 123.705 194.310 126.535 ;
        RECT 5.330 118.265 194.310 121.095 ;
        RECT 5.330 112.825 194.310 115.655 ;
        RECT 5.330 107.385 194.310 110.215 ;
        RECT 5.330 101.945 194.310 104.775 ;
        RECT 5.330 96.505 194.310 99.335 ;
        RECT 5.330 91.065 194.310 93.895 ;
        RECT 5.330 85.625 194.310 88.455 ;
        RECT 5.330 80.185 194.310 83.015 ;
        RECT 5.330 74.745 194.310 77.575 ;
        RECT 5.330 69.305 194.310 72.135 ;
        RECT 5.330 63.865 194.310 66.695 ;
        RECT 5.330 58.425 194.310 61.255 ;
        RECT 5.330 52.985 194.310 55.815 ;
        RECT 5.330 47.545 194.310 50.375 ;
        RECT 5.330 42.105 194.310 44.935 ;
        RECT 5.330 36.665 194.310 39.495 ;
        RECT 5.330 31.225 194.310 34.055 ;
        RECT 5.330 25.785 194.310 28.615 ;
        RECT 5.330 20.345 194.310 23.175 ;
        RECT 5.330 14.905 194.310 17.735 ;
        RECT 5.330 10.690 194.310 12.295 ;
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 5.520 4.800 194.120 187.920 ;
      LAYER met2 ;
        RECT 11.140 195.720 99.630 196.000 ;
        RECT 100.470 195.720 188.960 196.000 ;
        RECT 11.140 4.280 188.960 195.720 ;
        RECT 11.690 4.000 32.930 4.280 ;
        RECT 33.770 4.000 55.010 4.280 ;
        RECT 55.850 4.000 77.550 4.280 ;
        RECT 78.390 4.000 99.630 4.280 ;
        RECT 100.470 4.000 121.710 4.280 ;
        RECT 122.550 4.000 144.250 4.280 ;
        RECT 145.090 4.000 166.330 4.280 ;
        RECT 167.170 4.000 188.410 4.280 ;
      LAYER met3 ;
        RECT 21.040 10.715 176.240 187.845 ;
  END
END lfsr32
END LIBRARY

