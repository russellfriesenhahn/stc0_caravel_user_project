magic
tech sky130A
magscale 1 2
timestamp 1624325246
<< obsli1 >>
rect 1152 2647 244032 245105
<< obsm1 >>
rect 1152 2615 244032 245137
<< metal2 >>
rect 7604 247427 7660 248227
rect 22868 247427 22924 248227
rect 38228 247427 38284 248227
rect 53492 247427 53548 248227
rect 68852 247427 68908 248227
rect 84212 247427 84268 248227
rect 99476 247427 99532 248227
rect 114836 247427 114892 248227
rect 130196 247427 130252 248227
rect 145460 247427 145516 248227
rect 160820 247427 160876 248227
rect 176084 247427 176140 248227
rect 191444 247427 191500 248227
rect 206804 247427 206860 248227
rect 222068 247427 222124 248227
rect 237428 247427 237484 248227
<< obsm2 >>
rect 1556 247371 7548 247427
rect 7716 247371 22812 247427
rect 22980 247371 38172 247427
rect 38340 247371 53436 247427
rect 53604 247371 68796 247427
rect 68964 247371 84156 247427
rect 84324 247371 99420 247427
rect 99588 247371 114780 247427
rect 114948 247371 130140 247427
rect 130308 247371 145404 247427
rect 145572 247371 160764 247427
rect 160932 247371 176028 247427
rect 176196 247371 191388 247427
rect 191556 247371 206748 247427
rect 206916 247371 222012 247427
rect 222180 247371 237372 247427
rect 237540 247371 243530 247427
rect 1556 2616 243530 247371
<< metal3 >>
rect 0 241106 800 241226
rect 0 227342 800 227462
rect 244403 227342 245203 227462
rect 0 213578 800 213698
rect 0 199814 800 199934
rect 0 186050 800 186170
rect 244403 186050 245203 186170
rect 0 172286 800 172406
rect 0 158374 800 158494
rect 0 144610 800 144730
rect 244403 144610 245203 144730
rect 0 130846 800 130966
rect 0 117082 800 117202
rect 0 103318 800 103438
rect 244403 103318 245203 103438
rect 0 89554 800 89674
rect 0 75642 800 75762
rect 0 61878 800 61998
rect 244403 61878 245203 61998
rect 0 48114 800 48234
rect 0 34350 800 34470
rect 0 20586 800 20706
rect 244403 20586 245203 20706
rect 0 6822 800 6942
<< obsm3 >>
rect 800 241306 244403 245121
rect 880 241026 244403 241306
rect 800 227542 244403 241026
rect 880 227262 244323 227542
rect 800 213778 244403 227262
rect 880 213498 244403 213778
rect 800 200014 244403 213498
rect 880 199734 244403 200014
rect 800 186250 244403 199734
rect 880 185970 244323 186250
rect 800 172486 244403 185970
rect 880 172206 244403 172486
rect 800 158574 244403 172206
rect 880 158294 244403 158574
rect 800 144810 244403 158294
rect 880 144530 244323 144810
rect 800 131046 244403 144530
rect 880 130766 244403 131046
rect 800 117282 244403 130766
rect 880 117002 244403 117282
rect 800 103518 244403 117002
rect 880 103238 244323 103518
rect 800 89754 244403 103238
rect 880 89474 244403 89754
rect 800 75842 244403 89474
rect 880 75562 244403 75842
rect 800 62078 244403 75562
rect 880 61798 244323 62078
rect 800 48314 244403 61798
rect 880 48034 244403 48314
rect 800 34550 244403 48034
rect 880 34270 244403 34550
rect 800 20786 244403 34270
rect 880 20506 244323 20786
rect 800 7022 244403 20506
rect 880 6742 244403 7022
rect 800 2631 244403 6742
<< metal4 >>
rect 4256 2616 4576 245136
rect 4916 2664 5236 245088
rect 5576 2664 5896 245088
rect 6236 2664 6556 245088
rect 19616 2616 19936 245136
rect 20276 2664 20596 245088
rect 20936 2664 21256 245088
rect 21596 2664 21916 245088
rect 34976 2616 35296 245136
rect 35636 2664 35956 245088
rect 36296 2664 36616 245088
rect 36956 2664 37276 245088
rect 50336 2616 50656 245136
rect 50996 2664 51316 245088
rect 51656 2664 51976 245088
rect 52316 2664 52636 245088
rect 65696 2616 66016 245136
rect 66356 2664 66676 245088
rect 67016 2664 67336 245088
rect 67676 2664 67996 245088
rect 81056 2616 81376 245136
rect 81716 2664 82036 245088
rect 82376 2664 82696 245088
rect 83036 2664 83356 245088
rect 96416 2616 96736 245136
rect 97076 2664 97396 245088
rect 97736 2664 98056 245088
rect 98396 2664 98716 245088
rect 111776 2616 112096 245136
rect 112436 2664 112756 245088
rect 113096 2664 113416 245088
rect 113756 2664 114076 245088
rect 127136 2616 127456 245136
rect 127796 2664 128116 245088
rect 128456 2664 128776 245088
rect 129116 2664 129436 245088
rect 142496 2616 142816 245136
rect 143156 2664 143476 245088
rect 143816 2664 144136 245088
rect 144476 2664 144796 245088
rect 157856 2616 158176 245136
rect 158516 2664 158836 245088
rect 159176 2664 159496 245088
rect 159836 2664 160156 245088
rect 173216 2616 173536 245136
rect 173876 2664 174196 245088
rect 174536 2664 174856 245088
rect 175196 2664 175516 245088
rect 188576 2616 188896 245136
rect 189236 2664 189556 245088
rect 189896 2664 190216 245088
rect 190556 2664 190876 245088
rect 203936 2616 204256 245136
rect 204596 2664 204916 245088
rect 205256 2664 205576 245088
rect 205916 2664 206236 245088
rect 219296 2616 219616 245136
rect 219956 2664 220276 245088
rect 220616 2664 220936 245088
rect 221276 2664 221596 245088
rect 234656 2616 234976 245136
rect 235316 2664 235636 245088
rect 235976 2664 236296 245088
rect 236636 2664 236956 245088
<< obsm4 >>
rect 69759 7145 80976 204791
rect 81456 7145 81636 204791
rect 82116 7145 82296 204791
rect 82776 7145 82956 204791
rect 83436 7145 96336 204791
rect 96816 7145 96996 204791
rect 97476 7145 97656 204791
rect 98136 7145 98316 204791
rect 98796 7145 111696 204791
rect 112176 7145 112356 204791
rect 112836 7145 113016 204791
rect 113496 7145 113676 204791
rect 114156 7145 127056 204791
rect 127536 7145 127716 204791
rect 128196 7145 128376 204791
rect 128856 7145 129036 204791
rect 129516 7145 142416 204791
rect 142896 7145 143076 204791
rect 143556 7145 143736 204791
rect 144216 7145 144396 204791
rect 144876 7145 157776 204791
rect 158256 7145 158436 204791
rect 158916 7145 159096 204791
rect 159576 7145 159756 204791
rect 160236 7145 173136 204791
rect 173616 7145 173796 204791
rect 174276 7145 174456 204791
rect 174936 7145 175116 204791
rect 175596 7145 188496 204791
rect 188976 7145 189156 204791
rect 189636 7145 189816 204791
rect 190296 7145 190476 204791
rect 190956 7145 203856 204791
rect 204336 7145 204516 204791
rect 204996 7145 205176 204791
rect 205656 7145 205836 204791
rect 206316 7145 215937 204791
<< labels >>
rlabel metal3 s 0 48114 800 48234 6 ARstb
port 1 nsew signal input
rlabel metal3 s 0 20586 800 20706 6 ClkIngress
port 2 nsew signal input
rlabel metal3 s 244403 186050 245203 186170 6 ED[0]
port 3 nsew signal output
rlabel metal3 s 244403 103318 245203 103438 6 ED[1]
port 4 nsew signal output
rlabel metal3 s 244403 20586 245203 20706 6 ED[2]
port 5 nsew signal output
rlabel metal2 s 222068 247427 222124 248227 6 ED[3]
port 6 nsew signal output
rlabel metal2 s 160820 247427 160876 248227 6 ED[4]
port 7 nsew signal output
rlabel metal2 s 130196 247427 130252 248227 6 ED[5]
port 8 nsew signal output
rlabel metal2 s 99476 247427 99532 248227 6 ED[6]
port 9 nsew signal output
rlabel metal2 s 68852 247427 68908 248227 6 ED[7]
port 10 nsew signal output
rlabel metal2 s 191444 247427 191500 248227 6 EValid
port 11 nsew signal output
rlabel metal2 s 38228 247427 38284 248227 6 ID[0]
port 12 nsew signal input
rlabel metal2 s 7604 247427 7660 248227 6 ID[1]
port 13 nsew signal input
rlabel metal3 s 0 241106 800 241226 6 ID[2]
port 14 nsew signal input
rlabel metal3 s 0 213578 800 213698 6 ID[3]
port 15 nsew signal input
rlabel metal3 s 0 158374 800 158494 6 ID[4]
port 16 nsew signal input
rlabel metal3 s 0 130846 800 130966 6 ID[5]
port 17 nsew signal input
rlabel metal3 s 0 103318 800 103438 6 ID[6]
port 18 nsew signal input
rlabel metal3 s 0 75642 800 75762 6 ID[7]
port 19 nsew signal input
rlabel metal3 s 0 186050 800 186170 6 IValid
port 20 nsew signal input
rlabel metal3 s 244403 227342 245203 227462 6 io_oeb[0]
port 21 nsew signal output
rlabel metal2 s 22868 247427 22924 248227 6 io_oeb[10]
port 22 nsew signal output
rlabel metal3 s 0 227342 800 227462 6 io_oeb[11]
port 23 nsew signal output
rlabel metal3 s 0 199814 800 199934 6 io_oeb[12]
port 24 nsew signal output
rlabel metal3 s 0 172286 800 172406 6 io_oeb[13]
port 25 nsew signal output
rlabel metal3 s 0 144610 800 144730 6 io_oeb[14]
port 26 nsew signal output
rlabel metal3 s 0 117082 800 117202 6 io_oeb[15]
port 27 nsew signal output
rlabel metal3 s 0 89554 800 89674 6 io_oeb[16]
port 28 nsew signal output
rlabel metal3 s 0 61878 800 61998 6 io_oeb[17]
port 29 nsew signal output
rlabel metal3 s 0 34350 800 34470 6 io_oeb[18]
port 30 nsew signal output
rlabel metal3 s 0 6822 800 6942 6 io_oeb[19]
port 31 nsew signal output
rlabel metal3 s 244403 144610 245203 144730 6 io_oeb[1]
port 32 nsew signal output
rlabel metal3 s 244403 61878 245203 61998 6 io_oeb[2]
port 33 nsew signal output
rlabel metal2 s 237428 247427 237484 248227 6 io_oeb[3]
port 34 nsew signal output
rlabel metal2 s 206804 247427 206860 248227 6 io_oeb[4]
port 35 nsew signal output
rlabel metal2 s 176084 247427 176140 248227 6 io_oeb[5]
port 36 nsew signal output
rlabel metal2 s 145460 247427 145516 248227 6 io_oeb[6]
port 37 nsew signal output
rlabel metal2 s 114836 247427 114892 248227 6 io_oeb[7]
port 38 nsew signal output
rlabel metal2 s 84212 247427 84268 248227 6 io_oeb[8]
port 39 nsew signal output
rlabel metal2 s 53492 247427 53548 248227 6 io_oeb[9]
port 40 nsew signal output
rlabel metal4 s 219296 2616 219616 245136 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 188576 2616 188896 245136 6 vccd1
port 42 nsew power bidirectional
rlabel metal4 s 157856 2616 158176 245136 6 vccd1
port 43 nsew power bidirectional
rlabel metal4 s 127136 2616 127456 245136 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 96416 2616 96736 245136 6 vccd1
port 45 nsew power bidirectional
rlabel metal4 s 65696 2616 66016 245136 6 vccd1
port 46 nsew power bidirectional
rlabel metal4 s 34976 2616 35296 245136 6 vccd1
port 47 nsew power bidirectional
rlabel metal4 s 4256 2616 4576 245136 6 vccd1
port 48 nsew power bidirectional
rlabel metal4 s 234656 2616 234976 245136 6 vssd1
port 49 nsew ground bidirectional
rlabel metal4 s 203936 2616 204256 245136 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 173216 2616 173536 245136 6 vssd1
port 51 nsew ground bidirectional
rlabel metal4 s 142496 2616 142816 245136 6 vssd1
port 52 nsew ground bidirectional
rlabel metal4 s 111776 2616 112096 245136 6 vssd1
port 53 nsew ground bidirectional
rlabel metal4 s 81056 2616 81376 245136 6 vssd1
port 54 nsew ground bidirectional
rlabel metal4 s 50336 2616 50656 245136 6 vssd1
port 55 nsew ground bidirectional
rlabel metal4 s 19616 2616 19936 245136 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 219956 2664 220276 245088 6 vccd2
port 57 nsew power bidirectional
rlabel metal4 s 189236 2664 189556 245088 6 vccd2
port 58 nsew power bidirectional
rlabel metal4 s 158516 2664 158836 245088 6 vccd2
port 59 nsew power bidirectional
rlabel metal4 s 127796 2664 128116 245088 6 vccd2
port 60 nsew power bidirectional
rlabel metal4 s 97076 2664 97396 245088 6 vccd2
port 61 nsew power bidirectional
rlabel metal4 s 66356 2664 66676 245088 6 vccd2
port 62 nsew power bidirectional
rlabel metal4 s 35636 2664 35956 245088 6 vccd2
port 63 nsew power bidirectional
rlabel metal4 s 4916 2664 5236 245088 6 vccd2
port 64 nsew power bidirectional
rlabel metal4 s 235316 2664 235636 245088 6 vssd2
port 65 nsew ground bidirectional
rlabel metal4 s 204596 2664 204916 245088 6 vssd2
port 66 nsew ground bidirectional
rlabel metal4 s 173876 2664 174196 245088 6 vssd2
port 67 nsew ground bidirectional
rlabel metal4 s 143156 2664 143476 245088 6 vssd2
port 68 nsew ground bidirectional
rlabel metal4 s 112436 2664 112756 245088 6 vssd2
port 69 nsew ground bidirectional
rlabel metal4 s 81716 2664 82036 245088 6 vssd2
port 70 nsew ground bidirectional
rlabel metal4 s 50996 2664 51316 245088 6 vssd2
port 71 nsew ground bidirectional
rlabel metal4 s 20276 2664 20596 245088 6 vssd2
port 72 nsew ground bidirectional
rlabel metal4 s 220616 2664 220936 245088 6 vdda1
port 73 nsew power bidirectional
rlabel metal4 s 189896 2664 190216 245088 6 vdda1
port 74 nsew power bidirectional
rlabel metal4 s 159176 2664 159496 245088 6 vdda1
port 75 nsew power bidirectional
rlabel metal4 s 128456 2664 128776 245088 6 vdda1
port 76 nsew power bidirectional
rlabel metal4 s 97736 2664 98056 245088 6 vdda1
port 77 nsew power bidirectional
rlabel metal4 s 67016 2664 67336 245088 6 vdda1
port 78 nsew power bidirectional
rlabel metal4 s 36296 2664 36616 245088 6 vdda1
port 79 nsew power bidirectional
rlabel metal4 s 5576 2664 5896 245088 6 vdda1
port 80 nsew power bidirectional
rlabel metal4 s 235976 2664 236296 245088 6 vssa1
port 81 nsew ground bidirectional
rlabel metal4 s 205256 2664 205576 245088 6 vssa1
port 82 nsew ground bidirectional
rlabel metal4 s 174536 2664 174856 245088 6 vssa1
port 83 nsew ground bidirectional
rlabel metal4 s 143816 2664 144136 245088 6 vssa1
port 84 nsew ground bidirectional
rlabel metal4 s 113096 2664 113416 245088 6 vssa1
port 85 nsew ground bidirectional
rlabel metal4 s 82376 2664 82696 245088 6 vssa1
port 86 nsew ground bidirectional
rlabel metal4 s 51656 2664 51976 245088 6 vssa1
port 87 nsew ground bidirectional
rlabel metal4 s 20936 2664 21256 245088 6 vssa1
port 88 nsew ground bidirectional
rlabel metal4 s 221276 2664 221596 245088 6 vdda2
port 89 nsew power bidirectional
rlabel metal4 s 190556 2664 190876 245088 6 vdda2
port 90 nsew power bidirectional
rlabel metal4 s 159836 2664 160156 245088 6 vdda2
port 91 nsew power bidirectional
rlabel metal4 s 129116 2664 129436 245088 6 vdda2
port 92 nsew power bidirectional
rlabel metal4 s 98396 2664 98716 245088 6 vdda2
port 93 nsew power bidirectional
rlabel metal4 s 67676 2664 67996 245088 6 vdda2
port 94 nsew power bidirectional
rlabel metal4 s 36956 2664 37276 245088 6 vdda2
port 95 nsew power bidirectional
rlabel metal4 s 6236 2664 6556 245088 6 vdda2
port 96 nsew power bidirectional
rlabel metal4 s 236636 2664 236956 245088 6 vssa2
port 97 nsew ground bidirectional
rlabel metal4 s 205916 2664 206236 245088 6 vssa2
port 98 nsew ground bidirectional
rlabel metal4 s 175196 2664 175516 245088 6 vssa2
port 99 nsew ground bidirectional
rlabel metal4 s 144476 2664 144796 245088 6 vssa2
port 100 nsew ground bidirectional
rlabel metal4 s 113756 2664 114076 245088 6 vssa2
port 101 nsew ground bidirectional
rlabel metal4 s 83036 2664 83356 245088 6 vssa2
port 102 nsew ground bidirectional
rlabel metal4 s 52316 2664 52636 245088 6 vssa2
port 103 nsew ground bidirectional
rlabel metal4 s 21596 2664 21916 245088 6 vssa2
port 104 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 245203 248227
string LEFview TRUE
string GDS_FILE /project/openlane/stc0_core/runs/stc0_core/results/magic/stc0_core.gds
string GDS_END 80652818
string GDS_START 1526346
<< end >>

