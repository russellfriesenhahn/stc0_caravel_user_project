magic
tech sky130A
magscale 1 2
timestamp 1624324446
<< locali >>
rect 22937 8279 22971 8585
<< viali >>
rect 21097 37281 21131 37315
rect 20453 37213 20487 37247
rect 20453 36873 20487 36907
rect 20269 36669 20303 36703
rect 18705 21505 18739 21539
rect 19073 21437 19107 21471
rect 20499 21301 20533 21335
rect 19073 20961 19107 20995
rect 19993 20961 20027 20995
rect 20361 20961 20395 20995
rect 21787 20757 21821 20791
rect 19717 20417 19751 20451
rect 20085 20417 20119 20451
rect 21511 20213 21545 20247
rect 21649 19873 21683 19907
rect 22017 19805 22051 19839
rect 20223 19669 20257 19703
rect 20913 17697 20947 17731
rect 21281 17697 21315 17731
rect 22707 17493 22741 17527
rect 19993 14909 20027 14943
rect 20177 14773 20211 14807
rect 22753 14433 22787 14467
rect 22845 14229 22879 14263
rect 21925 12325 21959 12359
rect 20177 12257 20211 12291
rect 24133 12257 24167 12291
rect 25421 12257 25455 12291
rect 25237 12121 25271 12155
rect 19993 12053 20027 12087
rect 23397 12053 23431 12087
rect 24317 12053 24351 12087
rect 21649 11849 21683 11883
rect 23213 11781 23247 11815
rect 24041 11781 24075 11815
rect 21465 11645 21499 11679
rect 22753 11645 22787 11679
rect 23397 11645 23431 11679
rect 23857 11645 23891 11679
rect 24685 11645 24719 11679
rect 25329 11645 25363 11679
rect 22569 11509 22603 11543
rect 24501 11509 24535 11543
rect 25145 11509 25179 11543
rect 20729 11169 20763 11203
rect 23581 11169 23615 11203
rect 24225 11169 24259 11203
rect 25237 11169 25271 11203
rect 25881 11169 25915 11203
rect 22661 11101 22695 11135
rect 22937 11101 22971 11135
rect 21189 11033 21223 11067
rect 23397 11033 23431 11067
rect 24041 11033 24075 11067
rect 25421 11033 25455 11067
rect 26065 11033 26099 11067
rect 20545 10965 20579 10999
rect 22569 10761 22603 10795
rect 25605 10761 25639 10795
rect 20177 10693 20211 10727
rect 24041 10625 24075 10659
rect 19073 10557 19107 10591
rect 19717 10557 19751 10591
rect 20361 10557 20395 10591
rect 21005 10557 21039 10591
rect 21649 10557 21683 10591
rect 24317 10557 24351 10591
rect 24961 10557 24995 10591
rect 25421 10557 25455 10591
rect 26249 10557 26283 10591
rect 18889 10421 18923 10455
rect 19533 10421 19567 10455
rect 20821 10421 20855 10455
rect 21465 10421 21499 10455
rect 24777 10421 24811 10455
rect 26065 10421 26099 10455
rect 25881 10217 25915 10251
rect 19073 10081 19107 10115
rect 20361 10081 20395 10115
rect 21005 10081 21039 10115
rect 23673 10081 23707 10115
rect 25421 10081 25455 10115
rect 26065 10081 26099 10115
rect 26709 10081 26743 10115
rect 27353 10081 27387 10115
rect 27813 10081 27847 10115
rect 22937 10013 22971 10047
rect 23213 10013 23247 10047
rect 20821 9945 20855 9979
rect 26525 9945 26559 9979
rect 18889 9877 18923 9911
rect 20177 9877 20211 9911
rect 21465 9877 21499 9911
rect 23857 9877 23891 9911
rect 25237 9877 25271 9911
rect 27169 9877 27203 9911
rect 27997 9877 28031 9911
rect 19901 9537 19935 9571
rect 21649 9537 21683 9571
rect 22845 9537 22879 9571
rect 18613 9469 18647 9503
rect 19257 9469 19291 9503
rect 22569 9469 22603 9503
rect 26525 9469 26559 9503
rect 27997 9469 28031 9503
rect 28641 9469 28675 9503
rect 20177 9401 20211 9435
rect 26249 9401 26283 9435
rect 18797 9333 18831 9367
rect 19441 9333 19475 9367
rect 24317 9333 24351 9367
rect 24777 9333 24811 9367
rect 27813 9333 27847 9367
rect 28457 9333 28491 9367
rect 22017 9129 22051 9163
rect 28733 9129 28767 9163
rect 20545 9061 20579 9095
rect 25513 9061 25547 9095
rect 17601 8993 17635 9027
rect 18245 8993 18279 9027
rect 18889 8993 18923 9027
rect 25237 8993 25271 9027
rect 27629 8993 27663 9027
rect 28273 8993 28307 9027
rect 28917 8993 28951 9027
rect 20269 8925 20303 8959
rect 22477 8925 22511 8959
rect 22753 8925 22787 8959
rect 17785 8857 17819 8891
rect 19073 8857 19107 8891
rect 26985 8857 27019 8891
rect 28089 8857 28123 8891
rect 18429 8789 18463 8823
rect 24225 8789 24259 8823
rect 27445 8789 27479 8823
rect 19177 8585 19211 8619
rect 22937 8585 22971 8619
rect 25881 8585 25915 8619
rect 26525 8585 26559 8619
rect 19901 8449 19935 8483
rect 21649 8449 21683 8483
rect 19441 8381 19475 8415
rect 21373 8313 21407 8347
rect 24777 8449 24811 8483
rect 28089 8449 28123 8483
rect 23029 8381 23063 8415
rect 25237 8381 25271 8415
rect 26065 8381 26099 8415
rect 26709 8381 26743 8415
rect 27813 8381 27847 8415
rect 30205 8381 30239 8415
rect 23305 8313 23339 8347
rect 17693 8245 17727 8279
rect 22937 8245 22971 8279
rect 25421 8245 25455 8279
rect 29561 8245 29595 8279
rect 30021 8245 30055 8279
rect 19073 8041 19107 8075
rect 24317 8041 24351 8075
rect 27445 8041 27479 8075
rect 31125 8041 31159 8075
rect 17601 7973 17635 8007
rect 28917 7973 28951 8007
rect 16037 7905 16071 7939
rect 16865 7905 16899 7939
rect 17325 7905 17359 7939
rect 20361 7905 20395 7939
rect 29193 7905 29227 7939
rect 30665 7905 30699 7939
rect 31309 7905 31343 7939
rect 20637 7837 20671 7871
rect 22569 7837 22603 7871
rect 22845 7837 22879 7871
rect 25237 7837 25271 7871
rect 25513 7837 25547 7871
rect 26985 7837 27019 7871
rect 16221 7701 16255 7735
rect 16681 7701 16715 7735
rect 22109 7701 22143 7735
rect 30481 7701 30515 7735
rect 16405 7497 16439 7531
rect 22753 7497 22787 7531
rect 24961 7497 24995 7531
rect 31309 7497 31343 7531
rect 15117 7429 15151 7463
rect 30205 7429 30239 7463
rect 17693 7361 17727 7395
rect 17969 7361 18003 7395
rect 20177 7361 20211 7395
rect 24225 7361 24259 7395
rect 24501 7361 24535 7395
rect 26433 7361 26467 7395
rect 26709 7361 26743 7395
rect 28089 7361 28123 7395
rect 14933 7293 14967 7327
rect 15577 7293 15611 7327
rect 16221 7293 16255 7327
rect 19901 7293 19935 7327
rect 27813 7293 27847 7327
rect 30021 7293 30055 7327
rect 30849 7293 30883 7327
rect 31493 7293 31527 7327
rect 15761 7157 15795 7191
rect 19441 7157 19475 7191
rect 21649 7157 21683 7191
rect 29561 7157 29595 7191
rect 30665 7157 30699 7191
rect 20177 6953 20211 6987
rect 29193 6953 29227 6987
rect 30481 6953 30515 6987
rect 21649 6885 21683 6919
rect 27721 6885 27755 6919
rect 15117 6817 15151 6851
rect 21925 6817 21959 6851
rect 24133 6817 24167 6851
rect 26985 6817 27019 6851
rect 27445 6817 27479 6851
rect 30665 6817 30699 6851
rect 31125 6817 31159 6851
rect 31953 6817 31987 6851
rect 32597 6817 32631 6851
rect 15393 6749 15427 6783
rect 17325 6749 17359 6783
rect 17601 6749 17635 6783
rect 19073 6749 19107 6783
rect 23857 6749 23891 6783
rect 26709 6749 26743 6783
rect 22385 6681 22419 6715
rect 31769 6681 31803 6715
rect 16865 6613 16899 6647
rect 25237 6613 25271 6647
rect 31309 6613 31343 6647
rect 32413 6613 32447 6647
rect 14657 6409 14691 6443
rect 24317 6409 24351 6443
rect 30021 6409 30055 6443
rect 31309 6409 31343 6443
rect 14197 6341 14231 6375
rect 19441 6341 19475 6375
rect 16129 6273 16163 6307
rect 16405 6273 16439 6307
rect 17693 6273 17727 6307
rect 17969 6273 18003 6307
rect 21649 6273 21683 6307
rect 22845 6273 22879 6307
rect 14013 6205 14047 6239
rect 19901 6205 19935 6239
rect 22569 6205 22603 6239
rect 26525 6205 26559 6239
rect 27813 6205 27847 6239
rect 30205 6205 30239 6239
rect 30849 6205 30883 6239
rect 31493 6205 31527 6239
rect 32137 6205 32171 6239
rect 20177 6137 20211 6171
rect 26249 6137 26283 6171
rect 28089 6137 28123 6171
rect 24777 6069 24811 6103
rect 29561 6069 29595 6103
rect 30665 6069 30699 6103
rect 31953 6069 31987 6103
rect 13829 5865 13863 5899
rect 17325 5865 17359 5899
rect 24225 5865 24259 5899
rect 26985 5865 27019 5899
rect 22753 5797 22787 5831
rect 25513 5797 25547 5831
rect 13645 5729 13679 5763
rect 16865 5729 16899 5763
rect 19073 5729 19107 5763
rect 20269 5729 20303 5763
rect 22477 5729 22511 5763
rect 25237 5729 25271 5763
rect 29193 5729 29227 5763
rect 30665 5729 30699 5763
rect 31125 5729 31159 5763
rect 31953 5729 31987 5763
rect 32597 5729 32631 5763
rect 16589 5661 16623 5695
rect 18797 5661 18831 5695
rect 20545 5661 20579 5695
rect 28917 5661 28951 5695
rect 15117 5525 15151 5559
rect 22017 5525 22051 5559
rect 27445 5525 27479 5559
rect 30481 5525 30515 5559
rect 31309 5525 31343 5559
rect 31769 5525 31803 5559
rect 32413 5525 32447 5559
rect 17693 5321 17727 5355
rect 24869 5321 24903 5355
rect 30665 5321 30699 5355
rect 24409 5253 24443 5287
rect 31309 5253 31343 5287
rect 14105 5185 14139 5219
rect 19441 5185 19475 5219
rect 19901 5185 19935 5219
rect 20177 5185 20211 5219
rect 22661 5185 22695 5219
rect 22937 5185 22971 5219
rect 26617 5185 26651 5219
rect 14197 5117 14231 5151
rect 14657 5117 14691 5151
rect 29561 5117 29595 5151
rect 30205 5117 30239 5151
rect 30849 5117 30883 5151
rect 31493 5117 31527 5151
rect 14933 5049 14967 5083
rect 19165 5049 19199 5083
rect 26341 5049 26375 5083
rect 29285 5049 29319 5083
rect 16405 4981 16439 5015
rect 21649 4981 21683 5015
rect 27813 4981 27847 5015
rect 30021 4981 30055 5015
rect 15117 4777 15151 4811
rect 27905 4777 27939 4811
rect 22845 4709 22879 4743
rect 28457 4709 28491 4743
rect 16865 4641 16899 4675
rect 17325 4641 17359 4675
rect 22569 4641 22603 4675
rect 27077 4641 27111 4675
rect 28181 4641 28215 4675
rect 29193 4641 29227 4675
rect 30665 4641 30699 4675
rect 16589 4573 16623 4607
rect 21465 4573 21499 4607
rect 21833 4573 21867 4607
rect 24317 4573 24351 4607
rect 27445 4573 27479 4607
rect 28089 4573 28123 4607
rect 28549 4573 28583 4607
rect 19073 4505 19107 4539
rect 29009 4505 29043 4539
rect 17588 4437 17622 4471
rect 20039 4437 20073 4471
rect 25651 4437 25685 4471
rect 30481 4437 30515 4471
rect 16221 4233 16255 4267
rect 20164 4233 20198 4267
rect 25224 4233 25258 4267
rect 27813 4233 27847 4267
rect 17693 4097 17727 4131
rect 22661 4097 22695 4131
rect 28365 4097 28399 4131
rect 14933 4029 14967 4063
rect 15577 4029 15611 4063
rect 16405 4029 16439 4063
rect 19901 4029 19935 4063
rect 24409 4029 24443 4063
rect 24961 4029 24995 4063
rect 27997 4029 28031 4063
rect 28089 4029 28123 4063
rect 29101 4029 29135 4063
rect 29745 4029 29779 4063
rect 30205 4029 30239 4063
rect 17969 3961 18003 3995
rect 24133 3961 24167 3995
rect 28457 3961 28491 3995
rect 15117 3893 15151 3927
rect 15761 3893 15795 3927
rect 19441 3893 19475 3927
rect 21649 3893 21683 3927
rect 26709 3893 26743 3927
rect 28917 3893 28951 3927
rect 29561 3893 29595 3927
rect 30297 3893 30331 3927
rect 16865 3689 16899 3723
rect 19073 3689 19107 3723
rect 24317 3689 24351 3723
rect 26985 3689 27019 3723
rect 29377 3689 29411 3723
rect 17601 3621 17635 3655
rect 22845 3621 22879 3655
rect 25513 3621 25547 3655
rect 16037 3553 16071 3587
rect 16681 3553 16715 3587
rect 17325 3553 17359 3587
rect 22109 3553 22143 3587
rect 22569 3553 22603 3587
rect 25237 3553 25271 3587
rect 27445 3553 27479 3587
rect 28273 3553 28307 3587
rect 28917 3553 28951 3587
rect 29561 3553 29595 3587
rect 21833 3485 21867 3519
rect 27629 3417 27663 3451
rect 28089 3417 28123 3451
rect 16129 3349 16163 3383
rect 20361 3349 20395 3383
rect 28733 3349 28767 3383
rect 17877 3145 17911 3179
rect 18337 3145 18371 3179
rect 19441 3145 19475 3179
rect 19901 3145 19935 3179
rect 24317 3145 24351 3179
rect 26157 3145 26191 3179
rect 26617 3145 26651 3179
rect 25605 3077 25639 3111
rect 29101 3077 29135 3111
rect 30205 3077 30239 3111
rect 19257 3009 19291 3043
rect 21373 3009 21407 3043
rect 21649 3009 21683 3043
rect 22845 3009 22879 3043
rect 29745 3009 29779 3043
rect 17785 2941 17819 2975
rect 18061 2941 18095 2975
rect 18153 2941 18187 2975
rect 18797 2941 18831 2975
rect 18889 2941 18923 2975
rect 19165 2941 19199 2975
rect 22569 2941 22603 2975
rect 24777 2941 24811 2975
rect 25421 2941 25455 2975
rect 26341 2941 26375 2975
rect 26433 2941 26467 2975
rect 26709 2941 26743 2975
rect 27997 2941 28031 2975
rect 28641 2941 28675 2975
rect 30389 2941 30423 2975
rect 11161 2805 11195 2839
rect 24961 2805 24995 2839
rect 27813 2805 27847 2839
rect 28457 2805 28491 2839
rect 19349 2601 19383 2635
rect 22937 2601 22971 2635
rect 25605 2601 25639 2635
rect 26249 2601 26283 2635
rect 28365 2601 28399 2635
rect 11253 2533 11287 2567
rect 15761 2533 15795 2567
rect 18705 2533 18739 2567
rect 21741 2533 21775 2567
rect 33793 2533 33827 2567
rect 2421 2465 2455 2499
rect 2973 2465 3007 2499
rect 16681 2465 16715 2499
rect 18061 2465 18095 2499
rect 18797 2465 18831 2499
rect 19073 2465 19107 2499
rect 22017 2465 22051 2499
rect 24685 2465 24719 2499
rect 25789 2465 25823 2499
rect 26433 2465 26467 2499
rect 27077 2465 27111 2499
rect 28457 2465 28491 2499
rect 29101 2465 29135 2499
rect 29653 2465 29687 2499
rect 37289 2465 37323 2499
rect 37933 2465 37967 2499
rect 19165 2397 19199 2431
rect 20269 2397 20303 2431
rect 24409 2397 24443 2431
rect 2237 2329 2271 2363
rect 11069 2329 11103 2363
rect 15577 2329 15611 2363
rect 18245 2329 18279 2363
rect 28917 2329 28951 2363
rect 33609 2329 33643 2363
rect 37749 2329 37783 2363
rect 26893 2261 26927 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 38824 37562
rect 1104 37488 38824 37510
rect 20806 37272 20812 37324
rect 20864 37312 20870 37324
rect 21085 37315 21143 37321
rect 21085 37312 21097 37315
rect 20864 37284 21097 37312
rect 20864 37272 20870 37284
rect 21085 37281 21097 37284
rect 21131 37281 21143 37315
rect 21085 37275 21143 37281
rect 20438 37244 20444 37256
rect 20399 37216 20444 37244
rect 20438 37204 20444 37216
rect 20496 37204 20502 37256
rect 1104 37018 38824 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 38824 37018
rect 1104 36944 38824 36966
rect 20438 36904 20444 36916
rect 20399 36876 20444 36904
rect 20438 36864 20444 36876
rect 20496 36864 20502 36916
rect 19978 36660 19984 36712
rect 20036 36700 20042 36712
rect 20257 36703 20315 36709
rect 20257 36700 20269 36703
rect 20036 36672 20269 36700
rect 20036 36660 20042 36672
rect 20257 36669 20269 36672
rect 20303 36669 20315 36703
rect 20257 36663 20315 36669
rect 1104 36474 38824 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 38824 36474
rect 1104 36400 38824 36422
rect 1104 35930 38824 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 38824 35930
rect 1104 35856 38824 35878
rect 1104 35386 38824 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 38824 35386
rect 1104 35312 38824 35334
rect 1104 34842 38824 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 38824 34842
rect 1104 34768 38824 34790
rect 1104 34298 38824 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 38824 34298
rect 1104 34224 38824 34246
rect 1104 33754 38824 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 38824 33754
rect 1104 33680 38824 33702
rect 1104 33210 38824 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 38824 33210
rect 1104 33136 38824 33158
rect 1104 32666 38824 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 38824 32666
rect 1104 32592 38824 32614
rect 1104 32122 38824 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 38824 32122
rect 1104 32048 38824 32070
rect 1104 31578 38824 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 38824 31578
rect 1104 31504 38824 31526
rect 1104 31034 38824 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 38824 31034
rect 1104 30960 38824 30982
rect 1104 30490 38824 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 38824 30490
rect 1104 30416 38824 30438
rect 1104 29946 38824 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 38824 29946
rect 1104 29872 38824 29894
rect 1104 29402 38824 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 38824 29402
rect 1104 29328 38824 29350
rect 1104 28858 38824 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 38824 28858
rect 1104 28784 38824 28806
rect 1104 28314 38824 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 38824 28314
rect 1104 28240 38824 28262
rect 1104 27770 38824 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 38824 27770
rect 1104 27696 38824 27718
rect 1104 27226 38824 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 38824 27226
rect 1104 27152 38824 27174
rect 1104 26682 38824 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 38824 26682
rect 1104 26608 38824 26630
rect 1104 26138 38824 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 38824 26138
rect 1104 26064 38824 26086
rect 1104 25594 38824 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 38824 25594
rect 1104 25520 38824 25542
rect 1104 25050 38824 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 38824 25050
rect 1104 24976 38824 24998
rect 1104 24506 38824 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 38824 24506
rect 1104 24432 38824 24454
rect 1104 23962 38824 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 38824 23962
rect 1104 23888 38824 23910
rect 1104 23418 38824 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 38824 23418
rect 1104 23344 38824 23366
rect 1104 22874 38824 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 38824 22874
rect 1104 22800 38824 22822
rect 1104 22330 38824 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 38824 22330
rect 1104 22256 38824 22278
rect 1104 21786 38824 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 38824 21786
rect 1104 21712 38824 21734
rect 18693 21539 18751 21545
rect 18693 21505 18705 21539
rect 18739 21536 18751 21539
rect 19978 21536 19984 21548
rect 18739 21508 19984 21536
rect 18739 21505 18751 21508
rect 18693 21499 18751 21505
rect 19978 21496 19984 21508
rect 20036 21496 20042 21548
rect 19058 21468 19064 21480
rect 19019 21440 19064 21468
rect 19058 21428 19064 21440
rect 19116 21428 19122 21480
rect 20806 21400 20812 21412
rect 20102 21372 20812 21400
rect 20806 21360 20812 21372
rect 20864 21360 20870 21412
rect 20346 21292 20352 21344
rect 20404 21332 20410 21344
rect 20487 21335 20545 21341
rect 20487 21332 20499 21335
rect 20404 21304 20499 21332
rect 20404 21292 20410 21304
rect 20487 21301 20499 21304
rect 20533 21301 20545 21335
rect 20487 21295 20545 21301
rect 1104 21242 38824 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 38824 21242
rect 1104 21168 38824 21190
rect 20806 21088 20812 21140
rect 20864 21088 20870 21140
rect 20824 21046 20852 21088
rect 19058 20992 19064 21004
rect 19019 20964 19064 20992
rect 19058 20952 19064 20964
rect 19116 20952 19122 21004
rect 19978 20992 19984 21004
rect 19939 20964 19984 20992
rect 19978 20952 19984 20964
rect 20036 20952 20042 21004
rect 20346 20992 20352 21004
rect 20307 20964 20352 20992
rect 20346 20952 20352 20964
rect 20404 20952 20410 21004
rect 20898 20748 20904 20800
rect 20956 20788 20962 20800
rect 21775 20791 21833 20797
rect 21775 20788 21787 20791
rect 20956 20760 21787 20788
rect 20956 20748 20962 20760
rect 21775 20757 21787 20760
rect 21821 20757 21833 20791
rect 21775 20751 21833 20757
rect 1104 20698 38824 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 38824 20698
rect 1104 20624 38824 20646
rect 19705 20451 19763 20457
rect 19705 20417 19717 20451
rect 19751 20448 19763 20451
rect 19978 20448 19984 20460
rect 19751 20420 19984 20448
rect 19751 20417 19763 20420
rect 19705 20411 19763 20417
rect 19978 20408 19984 20420
rect 20036 20408 20042 20460
rect 20073 20451 20131 20457
rect 20073 20417 20085 20451
rect 20119 20448 20131 20451
rect 20898 20448 20904 20460
rect 20119 20420 20904 20448
rect 20119 20417 20131 20420
rect 20073 20411 20131 20417
rect 20898 20408 20904 20420
rect 20956 20408 20962 20460
rect 20806 20272 20812 20324
rect 20864 20272 20870 20324
rect 21499 20247 21557 20253
rect 21499 20213 21511 20247
rect 21545 20244 21557 20247
rect 21634 20244 21640 20256
rect 21545 20216 21640 20244
rect 21545 20213 21557 20216
rect 21499 20207 21557 20213
rect 21634 20204 21640 20216
rect 21692 20204 21698 20256
rect 1104 20154 38824 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 38824 20154
rect 1104 20080 38824 20102
rect 20806 19932 20812 19984
rect 20864 19932 20870 19984
rect 21634 19904 21640 19916
rect 21595 19876 21640 19904
rect 21634 19864 21640 19876
rect 21692 19864 21698 19916
rect 22005 19839 22063 19845
rect 22005 19805 22017 19839
rect 22051 19836 22063 19839
rect 22094 19836 22100 19848
rect 22051 19808 22100 19836
rect 22051 19805 22063 19808
rect 22005 19799 22063 19805
rect 22094 19796 22100 19808
rect 22152 19796 22158 19848
rect 20211 19703 20269 19709
rect 20211 19669 20223 19703
rect 20257 19700 20269 19703
rect 21266 19700 21272 19712
rect 20257 19672 21272 19700
rect 20257 19669 20269 19672
rect 20211 19663 20269 19669
rect 21266 19660 21272 19672
rect 21324 19660 21330 19712
rect 1104 19610 38824 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 38824 19610
rect 1104 19536 38824 19558
rect 1104 19066 38824 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 38824 19066
rect 1104 18992 38824 19014
rect 1104 18522 38824 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 38824 18522
rect 1104 18448 38824 18470
rect 1104 17978 38824 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 38824 17978
rect 1104 17904 38824 17926
rect 20806 17824 20812 17876
rect 20864 17864 20870 17876
rect 20864 17836 21680 17864
rect 20864 17824 20870 17836
rect 21652 17782 21680 17836
rect 19978 17688 19984 17740
rect 20036 17728 20042 17740
rect 20901 17731 20959 17737
rect 20901 17728 20913 17731
rect 20036 17700 20913 17728
rect 20036 17688 20042 17700
rect 20901 17697 20913 17700
rect 20947 17697 20959 17731
rect 21266 17728 21272 17740
rect 21227 17700 21272 17728
rect 20901 17691 20959 17697
rect 21266 17688 21272 17700
rect 21324 17688 21330 17740
rect 22738 17533 22744 17536
rect 22695 17527 22744 17533
rect 22695 17493 22707 17527
rect 22741 17493 22744 17527
rect 22695 17487 22744 17493
rect 22738 17484 22744 17487
rect 22796 17484 22802 17536
rect 1104 17434 38824 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 38824 17434
rect 1104 17360 38824 17382
rect 1104 16890 38824 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 38824 16890
rect 1104 16816 38824 16838
rect 1104 16346 38824 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 38824 16346
rect 1104 16272 38824 16294
rect 1104 15802 38824 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 38824 15802
rect 1104 15728 38824 15750
rect 1104 15258 38824 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 38824 15258
rect 1104 15184 38824 15206
rect 19978 14940 19984 14952
rect 19939 14912 19984 14940
rect 19978 14900 19984 14912
rect 20036 14900 20042 14952
rect 20070 14764 20076 14816
rect 20128 14804 20134 14816
rect 20165 14807 20223 14813
rect 20165 14804 20177 14807
rect 20128 14776 20177 14804
rect 20128 14764 20134 14776
rect 20165 14773 20177 14776
rect 20211 14804 20223 14807
rect 20254 14804 20260 14816
rect 20211 14776 20260 14804
rect 20211 14773 20223 14776
rect 20165 14767 20223 14773
rect 20254 14764 20260 14776
rect 20312 14764 20318 14816
rect 1104 14714 38824 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 38824 14714
rect 1104 14640 38824 14662
rect 22738 14464 22744 14476
rect 22699 14436 22744 14464
rect 22738 14424 22744 14436
rect 22796 14424 22802 14476
rect 22833 14263 22891 14269
rect 22833 14229 22845 14263
rect 22879 14260 22891 14263
rect 23658 14260 23664 14272
rect 22879 14232 23664 14260
rect 22879 14229 22891 14232
rect 22833 14223 22891 14229
rect 23658 14220 23664 14232
rect 23716 14220 23722 14272
rect 1104 14170 38824 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 38824 14170
rect 1104 14096 38824 14118
rect 1104 13626 38824 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 38824 13626
rect 1104 13552 38824 13574
rect 1104 13082 38824 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 38824 13082
rect 1104 13008 38824 13030
rect 1104 12538 38824 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 38824 12538
rect 1104 12464 38824 12486
rect 21913 12359 21971 12365
rect 21913 12356 21925 12359
rect 6886 12328 21925 12356
rect 6638 12248 6644 12300
rect 6696 12288 6702 12300
rect 6886 12288 6914 12328
rect 21913 12325 21925 12328
rect 21959 12325 21971 12359
rect 21913 12319 21971 12325
rect 20162 12288 20168 12300
rect 6696 12260 6914 12288
rect 20123 12260 20168 12288
rect 6696 12248 6702 12260
rect 20162 12248 20168 12260
rect 20220 12248 20226 12300
rect 23658 12248 23664 12300
rect 23716 12288 23722 12300
rect 24121 12291 24179 12297
rect 24121 12288 24133 12291
rect 23716 12260 24133 12288
rect 23716 12248 23722 12260
rect 24121 12257 24133 12260
rect 24167 12288 24179 12291
rect 24670 12288 24676 12300
rect 24167 12260 24676 12288
rect 24167 12257 24179 12260
rect 24121 12251 24179 12257
rect 24670 12248 24676 12260
rect 24728 12248 24734 12300
rect 25406 12288 25412 12300
rect 25367 12260 25412 12288
rect 25406 12248 25412 12260
rect 25464 12248 25470 12300
rect 23290 12112 23296 12164
rect 23348 12152 23354 12164
rect 25225 12155 25283 12161
rect 25225 12152 25237 12155
rect 23348 12124 25237 12152
rect 23348 12112 23354 12124
rect 25225 12121 25237 12124
rect 25271 12121 25283 12155
rect 25225 12115 25283 12121
rect 19426 12044 19432 12096
rect 19484 12084 19490 12096
rect 19978 12084 19984 12096
rect 19484 12056 19984 12084
rect 19484 12044 19490 12056
rect 19978 12044 19984 12056
rect 20036 12044 20042 12096
rect 23382 12084 23388 12096
rect 23343 12056 23388 12084
rect 23382 12044 23388 12056
rect 23440 12044 23446 12096
rect 24305 12087 24363 12093
rect 24305 12053 24317 12087
rect 24351 12084 24363 12087
rect 25406 12084 25412 12096
rect 24351 12056 25412 12084
rect 24351 12053 24363 12056
rect 24305 12047 24363 12053
rect 25406 12044 25412 12056
rect 25464 12044 25470 12096
rect 1104 11994 38824 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 38824 11994
rect 1104 11920 38824 11942
rect 21637 11883 21695 11889
rect 21637 11849 21649 11883
rect 21683 11880 21695 11883
rect 22094 11880 22100 11892
rect 21683 11852 22100 11880
rect 21683 11849 21695 11852
rect 21637 11843 21695 11849
rect 22094 11840 22100 11852
rect 22152 11840 22158 11892
rect 21542 11772 21548 11824
rect 21600 11812 21606 11824
rect 23201 11815 23259 11821
rect 23201 11812 23213 11815
rect 21600 11784 23213 11812
rect 21600 11772 21606 11784
rect 23201 11781 23213 11784
rect 23247 11781 23259 11815
rect 23201 11775 23259 11781
rect 24029 11815 24087 11821
rect 24029 11781 24041 11815
rect 24075 11812 24087 11815
rect 24075 11784 24716 11812
rect 24075 11781 24087 11784
rect 24029 11775 24087 11781
rect 20898 11636 20904 11688
rect 20956 11676 20962 11688
rect 21453 11679 21511 11685
rect 21453 11676 21465 11679
rect 20956 11648 21465 11676
rect 20956 11636 20962 11648
rect 21453 11645 21465 11648
rect 21499 11645 21511 11679
rect 21453 11639 21511 11645
rect 22370 11636 22376 11688
rect 22428 11676 22434 11688
rect 22741 11679 22799 11685
rect 22741 11676 22753 11679
rect 22428 11648 22753 11676
rect 22428 11636 22434 11648
rect 22741 11645 22753 11648
rect 22787 11645 22799 11679
rect 22741 11639 22799 11645
rect 23385 11679 23443 11685
rect 23385 11645 23397 11679
rect 23431 11676 23443 11679
rect 23658 11676 23664 11688
rect 23431 11648 23664 11676
rect 23431 11645 23443 11648
rect 23385 11639 23443 11645
rect 22462 11568 22468 11620
rect 22520 11608 22526 11620
rect 23400 11608 23428 11639
rect 23658 11636 23664 11648
rect 23716 11636 23722 11688
rect 24688 11685 24716 11784
rect 23845 11679 23903 11685
rect 23845 11645 23857 11679
rect 23891 11645 23903 11679
rect 23845 11639 23903 11645
rect 24673 11679 24731 11685
rect 24673 11645 24685 11679
rect 24719 11676 24731 11679
rect 25222 11676 25228 11688
rect 24719 11648 25228 11676
rect 24719 11645 24731 11648
rect 24673 11639 24731 11645
rect 22520 11580 23428 11608
rect 23860 11608 23888 11639
rect 25222 11636 25228 11648
rect 25280 11636 25286 11688
rect 25317 11679 25375 11685
rect 25317 11645 25329 11679
rect 25363 11676 25375 11679
rect 25406 11676 25412 11688
rect 25363 11648 25412 11676
rect 25363 11645 25375 11648
rect 25317 11639 25375 11645
rect 25406 11636 25412 11648
rect 25464 11676 25470 11688
rect 27982 11676 27988 11688
rect 25464 11648 27988 11676
rect 25464 11636 25470 11648
rect 27982 11636 27988 11648
rect 28040 11636 28046 11688
rect 25590 11608 25596 11620
rect 23860 11580 25596 11608
rect 22520 11568 22526 11580
rect 25590 11568 25596 11580
rect 25648 11568 25654 11620
rect 22557 11543 22615 11549
rect 22557 11509 22569 11543
rect 22603 11540 22615 11543
rect 23566 11540 23572 11552
rect 22603 11512 23572 11540
rect 22603 11509 22615 11512
rect 22557 11503 22615 11509
rect 23566 11500 23572 11512
rect 23624 11500 23630 11552
rect 24118 11500 24124 11552
rect 24176 11540 24182 11552
rect 24489 11543 24547 11549
rect 24489 11540 24501 11543
rect 24176 11512 24501 11540
rect 24176 11500 24182 11512
rect 24489 11509 24501 11512
rect 24535 11509 24547 11543
rect 24489 11503 24547 11509
rect 24578 11500 24584 11552
rect 24636 11540 24642 11552
rect 25133 11543 25191 11549
rect 25133 11540 25145 11543
rect 24636 11512 25145 11540
rect 24636 11500 24642 11512
rect 25133 11509 25145 11512
rect 25179 11509 25191 11543
rect 25133 11503 25191 11509
rect 1104 11450 38824 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 38824 11450
rect 1104 11376 38824 11398
rect 20732 11308 23428 11336
rect 20732 11209 20760 11308
rect 23400 11280 23428 11308
rect 20990 11228 20996 11280
rect 21048 11268 21054 11280
rect 21048 11240 21482 11268
rect 21048 11228 21054 11240
rect 23382 11228 23388 11280
rect 23440 11268 23446 11280
rect 23440 11240 25912 11268
rect 23440 11228 23446 11240
rect 20717 11203 20775 11209
rect 20717 11169 20729 11203
rect 20763 11169 20775 11203
rect 23566 11200 23572 11212
rect 23479 11172 23572 11200
rect 20717 11163 20775 11169
rect 23566 11160 23572 11172
rect 23624 11160 23630 11212
rect 23658 11160 23664 11212
rect 23716 11200 23722 11212
rect 24213 11203 24271 11209
rect 24213 11200 24225 11203
rect 23716 11172 24225 11200
rect 23716 11160 23722 11172
rect 24213 11169 24225 11172
rect 24259 11200 24271 11203
rect 25222 11200 25228 11212
rect 24259 11172 25084 11200
rect 25135 11172 25228 11200
rect 24259 11169 24271 11172
rect 24213 11163 24271 11169
rect 22646 11132 22652 11144
rect 22607 11104 22652 11132
rect 22646 11092 22652 11104
rect 22704 11092 22710 11144
rect 22925 11135 22983 11141
rect 22925 11101 22937 11135
rect 22971 11132 22983 11135
rect 23198 11132 23204 11144
rect 22971 11104 23204 11132
rect 22971 11101 22983 11104
rect 22925 11095 22983 11101
rect 23198 11092 23204 11104
rect 23256 11092 23262 11144
rect 23584 11132 23612 11160
rect 24762 11132 24768 11144
rect 23584 11104 24768 11132
rect 24762 11092 24768 11104
rect 24820 11092 24826 11144
rect 21174 11064 21180 11076
rect 21135 11036 21180 11064
rect 21174 11024 21180 11036
rect 21232 11024 21238 11076
rect 23385 11067 23443 11073
rect 23385 11064 23397 11067
rect 22848 11036 23397 11064
rect 19702 10956 19708 11008
rect 19760 10996 19766 11008
rect 20162 10996 20168 11008
rect 19760 10968 20168 10996
rect 19760 10956 19766 10968
rect 20162 10956 20168 10968
rect 20220 10996 20226 11008
rect 20533 10999 20591 11005
rect 20533 10996 20545 10999
rect 20220 10968 20545 10996
rect 20220 10956 20226 10968
rect 20533 10965 20545 10968
rect 20579 10965 20591 10999
rect 20533 10959 20591 10965
rect 22278 10956 22284 11008
rect 22336 10996 22342 11008
rect 22848 10996 22876 11036
rect 23385 11033 23397 11036
rect 23431 11033 23443 11067
rect 23385 11027 23443 11033
rect 23658 11024 23664 11076
rect 23716 11064 23722 11076
rect 24029 11067 24087 11073
rect 24029 11064 24041 11067
rect 23716 11036 24041 11064
rect 23716 11024 23722 11036
rect 24029 11033 24041 11036
rect 24075 11033 24087 11067
rect 24029 11027 24087 11033
rect 22336 10968 22876 10996
rect 22336 10956 22342 10968
rect 23198 10956 23204 11008
rect 23256 10996 23262 11008
rect 24394 10996 24400 11008
rect 23256 10968 24400 10996
rect 23256 10956 23262 10968
rect 24394 10956 24400 10968
rect 24452 10956 24458 11008
rect 25056 10996 25084 11172
rect 25222 11160 25228 11172
rect 25280 11160 25286 11212
rect 25884 11209 25912 11240
rect 25869 11203 25927 11209
rect 25869 11169 25881 11203
rect 25915 11169 25927 11203
rect 25869 11163 25927 11169
rect 25240 11132 25268 11160
rect 26234 11132 26240 11144
rect 25240 11104 26240 11132
rect 26234 11092 26240 11104
rect 26292 11092 26298 11144
rect 25409 11067 25467 11073
rect 25409 11033 25421 11067
rect 25455 11064 25467 11067
rect 25682 11064 25688 11076
rect 25455 11036 25688 11064
rect 25455 11033 25467 11036
rect 25409 11027 25467 11033
rect 25682 11024 25688 11036
rect 25740 11024 25746 11076
rect 25774 11024 25780 11076
rect 25832 11064 25838 11076
rect 26053 11067 26111 11073
rect 26053 11064 26065 11067
rect 25832 11036 26065 11064
rect 25832 11024 25838 11036
rect 26053 11033 26065 11036
rect 26099 11033 26111 11067
rect 26053 11027 26111 11033
rect 26142 10996 26148 11008
rect 25056 10968 26148 10996
rect 26142 10956 26148 10968
rect 26200 10956 26206 11008
rect 1104 10906 38824 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 38824 10906
rect 1104 10832 38824 10854
rect 22557 10795 22615 10801
rect 22557 10761 22569 10795
rect 22603 10792 22615 10795
rect 22646 10792 22652 10804
rect 22603 10764 22652 10792
rect 22603 10761 22615 10764
rect 22557 10755 22615 10761
rect 22646 10752 22652 10764
rect 22704 10752 22710 10804
rect 25590 10792 25596 10804
rect 25551 10764 25596 10792
rect 25590 10752 25596 10764
rect 25648 10792 25654 10804
rect 30006 10792 30012 10804
rect 25648 10764 30012 10792
rect 25648 10752 25654 10764
rect 30006 10752 30012 10764
rect 30064 10752 30070 10804
rect 19058 10684 19064 10736
rect 19116 10724 19122 10736
rect 20165 10727 20223 10733
rect 20165 10724 20177 10727
rect 19116 10696 20177 10724
rect 19116 10684 19122 10696
rect 20165 10693 20177 10696
rect 20211 10693 20223 10727
rect 20165 10687 20223 10693
rect 23566 10656 23572 10668
rect 20364 10628 23572 10656
rect 19061 10591 19119 10597
rect 19061 10557 19073 10591
rect 19107 10588 19119 10591
rect 19426 10588 19432 10600
rect 19107 10560 19432 10588
rect 19107 10557 19119 10560
rect 19061 10551 19119 10557
rect 19426 10548 19432 10560
rect 19484 10548 19490 10600
rect 19702 10588 19708 10600
rect 19663 10560 19708 10588
rect 19702 10548 19708 10560
rect 19760 10548 19766 10600
rect 19886 10548 19892 10600
rect 19944 10588 19950 10600
rect 20364 10597 20392 10628
rect 23566 10616 23572 10628
rect 23624 10616 23630 10668
rect 24029 10659 24087 10665
rect 24029 10625 24041 10659
rect 24075 10656 24087 10659
rect 27062 10656 27068 10668
rect 24075 10628 27068 10656
rect 24075 10625 24087 10628
rect 24029 10619 24087 10625
rect 27062 10616 27068 10628
rect 27120 10616 27126 10668
rect 20349 10591 20407 10597
rect 20349 10588 20361 10591
rect 19944 10560 20361 10588
rect 19944 10548 19950 10560
rect 20349 10557 20361 10560
rect 20395 10557 20407 10591
rect 20349 10551 20407 10557
rect 20806 10548 20812 10600
rect 20864 10588 20870 10600
rect 20993 10591 21051 10597
rect 20993 10588 21005 10591
rect 20864 10560 21005 10588
rect 20864 10548 20870 10560
rect 20993 10557 21005 10560
rect 21039 10588 21051 10591
rect 21637 10591 21695 10597
rect 21637 10588 21649 10591
rect 21039 10560 21649 10588
rect 21039 10557 21051 10560
rect 20993 10551 21051 10557
rect 21637 10557 21649 10560
rect 21683 10588 21695 10591
rect 22370 10588 22376 10600
rect 21683 10560 22376 10588
rect 21683 10557 21695 10560
rect 21637 10551 21695 10557
rect 22370 10548 22376 10560
rect 22428 10548 22434 10600
rect 24305 10591 24363 10597
rect 24305 10557 24317 10591
rect 24351 10588 24363 10591
rect 24394 10588 24400 10600
rect 24351 10560 24400 10588
rect 24351 10557 24363 10560
rect 24305 10551 24363 10557
rect 24394 10548 24400 10560
rect 24452 10548 24458 10600
rect 24762 10548 24768 10600
rect 24820 10588 24826 10600
rect 24949 10591 25007 10597
rect 24949 10588 24961 10591
rect 24820 10560 24961 10588
rect 24820 10548 24826 10560
rect 24949 10557 24961 10560
rect 24995 10557 25007 10591
rect 24949 10551 25007 10557
rect 25409 10591 25467 10597
rect 25409 10557 25421 10591
rect 25455 10557 25467 10591
rect 26234 10588 26240 10600
rect 26195 10560 26240 10588
rect 25409 10551 25467 10557
rect 22646 10480 22652 10532
rect 22704 10520 22710 10532
rect 22704 10492 22862 10520
rect 22704 10480 22710 10492
rect 24670 10480 24676 10532
rect 24728 10520 24734 10532
rect 25424 10520 25452 10551
rect 26234 10548 26240 10560
rect 26292 10548 26298 10600
rect 24728 10492 25452 10520
rect 24728 10480 24734 10492
rect 18877 10455 18935 10461
rect 18877 10421 18889 10455
rect 18923 10452 18935 10455
rect 19242 10452 19248 10464
rect 18923 10424 19248 10452
rect 18923 10421 18935 10424
rect 18877 10415 18935 10421
rect 19242 10412 19248 10424
rect 19300 10412 19306 10464
rect 19334 10412 19340 10464
rect 19392 10452 19398 10464
rect 19521 10455 19579 10461
rect 19521 10452 19533 10455
rect 19392 10424 19533 10452
rect 19392 10412 19398 10424
rect 19521 10421 19533 10424
rect 19567 10421 19579 10455
rect 19521 10415 19579 10421
rect 20346 10412 20352 10464
rect 20404 10452 20410 10464
rect 20809 10455 20867 10461
rect 20809 10452 20821 10455
rect 20404 10424 20821 10452
rect 20404 10412 20410 10424
rect 20809 10421 20821 10424
rect 20855 10421 20867 10455
rect 20809 10415 20867 10421
rect 21266 10412 21272 10464
rect 21324 10452 21330 10464
rect 21453 10455 21511 10461
rect 21453 10452 21465 10455
rect 21324 10424 21465 10452
rect 21324 10412 21330 10424
rect 21453 10421 21465 10424
rect 21499 10421 21511 10455
rect 21453 10415 21511 10421
rect 22738 10412 22744 10464
rect 22796 10452 22802 10464
rect 24765 10455 24823 10461
rect 24765 10452 24777 10455
rect 22796 10424 24777 10452
rect 22796 10412 22802 10424
rect 24765 10421 24777 10424
rect 24811 10421 24823 10455
rect 24765 10415 24823 10421
rect 25958 10412 25964 10464
rect 26016 10452 26022 10464
rect 26053 10455 26111 10461
rect 26053 10452 26065 10455
rect 26016 10424 26065 10452
rect 26016 10412 26022 10424
rect 26053 10421 26065 10424
rect 26099 10421 26111 10455
rect 26053 10415 26111 10421
rect 1104 10362 38824 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 38824 10362
rect 1104 10288 38824 10310
rect 25774 10248 25780 10260
rect 19076 10220 25780 10248
rect 19076 10121 19104 10220
rect 25774 10208 25780 10220
rect 25832 10208 25838 10260
rect 25869 10251 25927 10257
rect 25869 10217 25881 10251
rect 25915 10217 25927 10251
rect 25869 10211 25927 10217
rect 19242 10140 19248 10192
rect 19300 10180 19306 10192
rect 19426 10180 19432 10192
rect 19300 10152 19432 10180
rect 19300 10140 19306 10152
rect 19426 10140 19432 10152
rect 19484 10140 19490 10192
rect 25884 10180 25912 10211
rect 22494 10152 25912 10180
rect 19061 10115 19119 10121
rect 19061 10081 19073 10115
rect 19107 10081 19119 10115
rect 19061 10075 19119 10081
rect 19794 10072 19800 10124
rect 19852 10112 19858 10124
rect 20346 10112 20352 10124
rect 19852 10084 20352 10112
rect 19852 10072 19858 10084
rect 20346 10072 20352 10084
rect 20404 10072 20410 10124
rect 20993 10115 21051 10121
rect 20993 10081 21005 10115
rect 21039 10081 21051 10115
rect 23661 10115 23719 10121
rect 23661 10112 23673 10115
rect 20993 10075 21051 10081
rect 23584 10084 23673 10112
rect 20898 10044 20904 10056
rect 18892 10016 20904 10044
rect 18506 9868 18512 9920
rect 18564 9908 18570 9920
rect 18892 9917 18920 10016
rect 20898 10004 20904 10016
rect 20956 10004 20962 10056
rect 20806 9976 20812 9988
rect 20767 9948 20812 9976
rect 20806 9936 20812 9948
rect 20864 9936 20870 9988
rect 21008 9976 21036 10075
rect 22922 10044 22928 10056
rect 22883 10016 22928 10044
rect 22922 10004 22928 10016
rect 22980 10004 22986 10056
rect 23198 10044 23204 10056
rect 23159 10016 23204 10044
rect 23198 10004 23204 10016
rect 23256 10004 23262 10056
rect 21008 9948 21588 9976
rect 18877 9911 18935 9917
rect 18877 9908 18889 9911
rect 18564 9880 18889 9908
rect 18564 9868 18570 9880
rect 18877 9877 18889 9880
rect 18923 9877 18935 9911
rect 18877 9871 18935 9877
rect 19242 9868 19248 9920
rect 19300 9908 19306 9920
rect 20165 9911 20223 9917
rect 20165 9908 20177 9911
rect 19300 9880 20177 9908
rect 19300 9868 19306 9880
rect 20165 9877 20177 9880
rect 20211 9877 20223 9911
rect 20165 9871 20223 9877
rect 20714 9868 20720 9920
rect 20772 9908 20778 9920
rect 21453 9911 21511 9917
rect 21453 9908 21465 9911
rect 20772 9880 21465 9908
rect 20772 9868 20778 9880
rect 21453 9877 21465 9880
rect 21499 9877 21511 9911
rect 21560 9908 21588 9948
rect 23584 9908 23612 10084
rect 23661 10081 23673 10084
rect 23707 10112 23719 10115
rect 24670 10112 24676 10124
rect 23707 10084 24676 10112
rect 23707 10081 23719 10084
rect 23661 10075 23719 10081
rect 24670 10072 24676 10084
rect 24728 10072 24734 10124
rect 24762 10072 24768 10124
rect 24820 10112 24826 10124
rect 25409 10115 25467 10121
rect 25409 10112 25421 10115
rect 24820 10084 25421 10112
rect 24820 10072 24826 10084
rect 25409 10081 25421 10084
rect 25455 10081 25467 10115
rect 25409 10075 25467 10081
rect 26053 10115 26111 10121
rect 26053 10081 26065 10115
rect 26099 10112 26111 10115
rect 26142 10112 26148 10124
rect 26099 10084 26148 10112
rect 26099 10081 26111 10084
rect 26053 10075 26111 10081
rect 26142 10072 26148 10084
rect 26200 10072 26206 10124
rect 26234 10072 26240 10124
rect 26292 10112 26298 10124
rect 26697 10115 26755 10121
rect 26697 10112 26709 10115
rect 26292 10084 26709 10112
rect 26292 10072 26298 10084
rect 26697 10081 26709 10084
rect 26743 10112 26755 10115
rect 27154 10112 27160 10124
rect 26743 10084 27160 10112
rect 26743 10081 26755 10084
rect 26697 10075 26755 10081
rect 27154 10072 27160 10084
rect 27212 10072 27218 10124
rect 27338 10112 27344 10124
rect 27299 10084 27344 10112
rect 27338 10072 27344 10084
rect 27396 10072 27402 10124
rect 27801 10115 27859 10121
rect 27801 10081 27813 10115
rect 27847 10081 27859 10115
rect 27801 10075 27859 10081
rect 25222 10044 25228 10056
rect 21560 9880 23612 9908
rect 23676 10016 25228 10044
rect 23676 9908 23704 10016
rect 25222 10004 25228 10016
rect 25280 10004 25286 10056
rect 25774 10004 25780 10056
rect 25832 10044 25838 10056
rect 27816 10044 27844 10075
rect 25832 10016 27844 10044
rect 25832 10004 25838 10016
rect 23750 9936 23756 9988
rect 23808 9976 23814 9988
rect 26513 9979 26571 9985
rect 26513 9976 26525 9979
rect 23808 9948 26525 9976
rect 23808 9936 23814 9948
rect 26513 9945 26525 9948
rect 26559 9945 26571 9979
rect 26513 9939 26571 9945
rect 23845 9911 23903 9917
rect 23845 9908 23857 9911
rect 23676 9880 23857 9908
rect 21453 9871 21511 9877
rect 23845 9877 23857 9880
rect 23891 9877 23903 9911
rect 23845 9871 23903 9877
rect 24854 9868 24860 9920
rect 24912 9908 24918 9920
rect 25225 9911 25283 9917
rect 25225 9908 25237 9911
rect 24912 9880 25237 9908
rect 24912 9868 24918 9880
rect 25225 9877 25237 9880
rect 25271 9877 25283 9911
rect 27154 9908 27160 9920
rect 27115 9880 27160 9908
rect 25225 9871 25283 9877
rect 27154 9868 27160 9880
rect 27212 9868 27218 9920
rect 27985 9911 28043 9917
rect 27985 9877 27997 9911
rect 28031 9908 28043 9911
rect 31294 9908 31300 9920
rect 28031 9880 31300 9908
rect 28031 9877 28043 9880
rect 27985 9871 28043 9877
rect 31294 9868 31300 9880
rect 31352 9868 31358 9920
rect 1104 9818 38824 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 38824 9818
rect 1104 9744 38824 9766
rect 22664 9676 23888 9704
rect 22462 9636 22468 9648
rect 21192 9608 22468 9636
rect 17862 9528 17868 9580
rect 17920 9568 17926 9580
rect 19794 9568 19800 9580
rect 17920 9540 19800 9568
rect 17920 9528 17926 9540
rect 19260 9509 19288 9540
rect 19794 9528 19800 9540
rect 19852 9528 19858 9580
rect 19889 9571 19947 9577
rect 19889 9537 19901 9571
rect 19935 9568 19947 9571
rect 20254 9568 20260 9580
rect 19935 9540 20260 9568
rect 19935 9537 19947 9540
rect 19889 9531 19947 9537
rect 20254 9528 20260 9540
rect 20312 9528 20318 9580
rect 20622 9528 20628 9580
rect 20680 9568 20686 9580
rect 21192 9568 21220 9608
rect 22462 9596 22468 9608
rect 22520 9596 22526 9648
rect 20680 9540 21220 9568
rect 21637 9571 21695 9577
rect 20680 9528 20686 9540
rect 21637 9537 21649 9571
rect 21683 9568 21695 9571
rect 22664 9568 22692 9676
rect 23860 9636 23888 9676
rect 25240 9676 26464 9704
rect 25240 9636 25268 9676
rect 23860 9608 25268 9636
rect 26436 9636 26464 9676
rect 27798 9636 27804 9648
rect 26436 9608 27804 9636
rect 27798 9596 27804 9608
rect 27856 9596 27862 9648
rect 21683 9540 22692 9568
rect 22833 9571 22891 9577
rect 21683 9537 21695 9540
rect 21637 9531 21695 9537
rect 22833 9537 22845 9571
rect 22879 9568 22891 9571
rect 24302 9568 24308 9580
rect 22879 9540 24308 9568
rect 22879 9537 22891 9540
rect 22833 9531 22891 9537
rect 24302 9528 24308 9540
rect 24360 9528 24366 9580
rect 25222 9528 25228 9580
rect 25280 9568 25286 9580
rect 27338 9568 27344 9580
rect 25280 9540 27344 9568
rect 25280 9528 25286 9540
rect 27338 9528 27344 9540
rect 27396 9568 27402 9580
rect 27396 9540 28672 9568
rect 27396 9528 27402 9540
rect 18601 9503 18659 9509
rect 18601 9469 18613 9503
rect 18647 9469 18659 9503
rect 18601 9463 18659 9469
rect 19245 9503 19303 9509
rect 19245 9469 19257 9503
rect 19291 9469 19303 9503
rect 19245 9463 19303 9469
rect 18616 9432 18644 9463
rect 22094 9460 22100 9512
rect 22152 9500 22158 9512
rect 22554 9500 22560 9512
rect 22152 9472 22560 9500
rect 22152 9460 22158 9472
rect 22554 9460 22560 9472
rect 22612 9460 22618 9512
rect 26510 9460 26516 9512
rect 26568 9500 26574 9512
rect 27982 9500 27988 9512
rect 26568 9472 26613 9500
rect 27895 9472 27988 9500
rect 26568 9460 26574 9472
rect 27982 9460 27988 9472
rect 28040 9460 28046 9512
rect 28644 9509 28672 9540
rect 28629 9503 28687 9509
rect 28629 9469 28641 9503
rect 28675 9500 28687 9503
rect 30374 9500 30380 9512
rect 28675 9472 30380 9500
rect 28675 9469 28687 9472
rect 28629 9463 28687 9469
rect 30374 9460 30380 9472
rect 30432 9460 30438 9512
rect 19886 9432 19892 9444
rect 18616 9404 19892 9432
rect 19886 9392 19892 9404
rect 19944 9392 19950 9444
rect 20162 9432 20168 9444
rect 20123 9404 20168 9432
rect 20162 9392 20168 9404
rect 20220 9392 20226 9444
rect 22738 9432 22744 9444
rect 21390 9404 22744 9432
rect 22738 9392 22744 9404
rect 22796 9392 22802 9444
rect 24946 9432 24952 9444
rect 24058 9404 24952 9432
rect 24946 9392 24952 9404
rect 25004 9392 25010 9444
rect 25774 9392 25780 9444
rect 25832 9392 25838 9444
rect 26234 9432 26240 9444
rect 26195 9404 26240 9432
rect 26234 9392 26240 9404
rect 26292 9392 26298 9444
rect 28000 9432 28028 9460
rect 28902 9432 28908 9444
rect 28000 9404 28908 9432
rect 28902 9392 28908 9404
rect 28960 9392 28966 9444
rect 18690 9324 18696 9376
rect 18748 9364 18754 9376
rect 18785 9367 18843 9373
rect 18785 9364 18797 9367
rect 18748 9336 18797 9364
rect 18748 9324 18754 9336
rect 18785 9333 18797 9336
rect 18831 9333 18843 9367
rect 18785 9327 18843 9333
rect 19429 9367 19487 9373
rect 19429 9333 19441 9367
rect 19475 9364 19487 9367
rect 21082 9364 21088 9376
rect 19475 9336 21088 9364
rect 19475 9333 19487 9336
rect 19429 9327 19487 9333
rect 21082 9324 21088 9336
rect 21140 9324 21146 9376
rect 21726 9324 21732 9376
rect 21784 9364 21790 9376
rect 22646 9364 22652 9376
rect 21784 9336 22652 9364
rect 21784 9324 21790 9336
rect 22646 9324 22652 9336
rect 22704 9324 22710 9376
rect 23842 9324 23848 9376
rect 23900 9364 23906 9376
rect 24305 9367 24363 9373
rect 24305 9364 24317 9367
rect 23900 9336 24317 9364
rect 23900 9324 23906 9336
rect 24305 9333 24317 9336
rect 24351 9333 24363 9367
rect 24305 9327 24363 9333
rect 24765 9367 24823 9373
rect 24765 9333 24777 9367
rect 24811 9364 24823 9367
rect 25498 9364 25504 9376
rect 24811 9336 25504 9364
rect 24811 9333 24823 9336
rect 24765 9327 24823 9333
rect 25498 9324 25504 9336
rect 25556 9324 25562 9376
rect 25590 9324 25596 9376
rect 25648 9364 25654 9376
rect 27801 9367 27859 9373
rect 27801 9364 27813 9367
rect 25648 9336 27813 9364
rect 25648 9324 25654 9336
rect 27801 9333 27813 9336
rect 27847 9333 27859 9367
rect 28442 9364 28448 9376
rect 28403 9336 28448 9364
rect 27801 9327 27859 9333
rect 28442 9324 28448 9336
rect 28500 9324 28506 9376
rect 1104 9274 38824 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 38824 9274
rect 1104 9200 38824 9222
rect 22005 9163 22063 9169
rect 17604 9132 21956 9160
rect 17604 9033 17632 9132
rect 19978 9052 19984 9104
rect 20036 9092 20042 9104
rect 20533 9095 20591 9101
rect 20533 9092 20545 9095
rect 20036 9064 20545 9092
rect 20036 9052 20042 9064
rect 20533 9061 20545 9064
rect 20579 9061 20591 9095
rect 20533 9055 20591 9061
rect 21542 9052 21548 9104
rect 21600 9052 21606 9104
rect 21928 9092 21956 9132
rect 22005 9129 22017 9163
rect 22051 9160 22063 9163
rect 22922 9160 22928 9172
rect 22051 9132 22928 9160
rect 22051 9129 22063 9132
rect 22005 9123 22063 9129
rect 22922 9120 22928 9132
rect 22980 9120 22986 9172
rect 24670 9160 24676 9172
rect 23032 9132 24676 9160
rect 22370 9092 22376 9104
rect 21928 9064 22376 9092
rect 22370 9052 22376 9064
rect 22428 9092 22434 9104
rect 23032 9092 23060 9132
rect 24670 9120 24676 9132
rect 24728 9120 24734 9172
rect 24946 9120 24952 9172
rect 25004 9160 25010 9172
rect 28721 9163 28779 9169
rect 28721 9160 28733 9163
rect 25004 9132 28733 9160
rect 25004 9120 25010 9132
rect 28721 9129 28733 9132
rect 28767 9129 28779 9163
rect 28721 9123 28779 9129
rect 24578 9092 24584 9104
rect 22428 9064 23060 9092
rect 23966 9064 24584 9092
rect 22428 9052 22434 9064
rect 24578 9052 24584 9064
rect 24636 9052 24642 9104
rect 25498 9092 25504 9104
rect 25459 9064 25504 9092
rect 25498 9052 25504 9064
rect 25556 9052 25562 9104
rect 26510 9052 26516 9104
rect 26568 9052 26574 9104
rect 30466 9092 30472 9104
rect 27632 9064 30472 9092
rect 27632 9036 27660 9064
rect 30466 9052 30472 9064
rect 30524 9052 30530 9104
rect 17589 9027 17647 9033
rect 17589 8993 17601 9027
rect 17635 8993 17647 9027
rect 17589 8987 17647 8993
rect 17862 8984 17868 9036
rect 17920 9024 17926 9036
rect 18233 9027 18291 9033
rect 18233 9024 18245 9027
rect 17920 8996 18245 9024
rect 17920 8984 17926 8996
rect 18233 8993 18245 8996
rect 18279 8993 18291 9027
rect 18233 8987 18291 8993
rect 18877 9027 18935 9033
rect 18877 8993 18889 9027
rect 18923 9024 18935 9027
rect 20070 9024 20076 9036
rect 18923 8996 20076 9024
rect 18923 8993 18935 8996
rect 18877 8987 18935 8993
rect 17218 8916 17224 8968
rect 17276 8956 17282 8968
rect 18892 8956 18920 8987
rect 20070 8984 20076 8996
rect 20128 8984 20134 9036
rect 25130 8984 25136 9036
rect 25188 9024 25194 9036
rect 25225 9027 25283 9033
rect 25225 9024 25237 9027
rect 25188 8996 25237 9024
rect 25188 8984 25194 8996
rect 25225 8993 25237 8996
rect 25271 8993 25283 9027
rect 27614 9024 27620 9036
rect 27575 8996 27620 9024
rect 25225 8987 25283 8993
rect 27614 8984 27620 8996
rect 27672 8984 27678 9036
rect 28261 9027 28319 9033
rect 28261 8993 28273 9027
rect 28307 8993 28319 9027
rect 28902 9024 28908 9036
rect 28863 8996 28908 9024
rect 28261 8987 28319 8993
rect 17276 8928 18920 8956
rect 17276 8916 17282 8928
rect 19426 8916 19432 8968
rect 19484 8956 19490 8968
rect 20257 8959 20315 8965
rect 20257 8956 20269 8959
rect 19484 8928 20269 8956
rect 19484 8916 19490 8928
rect 20257 8925 20269 8928
rect 20303 8925 20315 8959
rect 21726 8956 21732 8968
rect 20257 8919 20315 8925
rect 20364 8928 21732 8956
rect 17773 8891 17831 8897
rect 17773 8857 17785 8891
rect 17819 8888 17831 8891
rect 19061 8891 19119 8897
rect 17819 8860 19012 8888
rect 17819 8857 17831 8860
rect 17773 8851 17831 8857
rect 18322 8780 18328 8832
rect 18380 8820 18386 8832
rect 18417 8823 18475 8829
rect 18417 8820 18429 8823
rect 18380 8792 18429 8820
rect 18380 8780 18386 8792
rect 18417 8789 18429 8792
rect 18463 8789 18475 8823
rect 18984 8820 19012 8860
rect 19061 8857 19073 8891
rect 19107 8888 19119 8891
rect 20364 8888 20392 8928
rect 21726 8916 21732 8928
rect 21784 8916 21790 8968
rect 22462 8956 22468 8968
rect 22423 8928 22468 8956
rect 22462 8916 22468 8928
rect 22520 8916 22526 8968
rect 22738 8956 22744 8968
rect 22699 8928 22744 8956
rect 22738 8916 22744 8928
rect 22796 8916 22802 8968
rect 28276 8956 28304 8987
rect 28902 8984 28908 8996
rect 28960 8984 28966 9036
rect 30190 8956 30196 8968
rect 25227 8928 28120 8956
rect 28276 8928 30196 8956
rect 25227 8888 25255 8928
rect 19107 8860 20392 8888
rect 24044 8860 25255 8888
rect 26973 8891 27031 8897
rect 19107 8857 19119 8860
rect 19061 8851 19119 8857
rect 20622 8820 20628 8832
rect 18984 8792 20628 8820
rect 18417 8783 18475 8789
rect 20622 8780 20628 8792
rect 20680 8780 20686 8832
rect 20898 8780 20904 8832
rect 20956 8820 20962 8832
rect 24044 8820 24072 8860
rect 26973 8857 26985 8891
rect 27019 8888 27031 8891
rect 27706 8888 27712 8900
rect 27019 8860 27712 8888
rect 27019 8857 27031 8860
rect 26973 8851 27031 8857
rect 27706 8848 27712 8860
rect 27764 8848 27770 8900
rect 28092 8897 28120 8928
rect 30190 8916 30196 8928
rect 30248 8916 30254 8968
rect 28077 8891 28135 8897
rect 28077 8857 28089 8891
rect 28123 8857 28135 8891
rect 28077 8851 28135 8857
rect 24210 8820 24216 8832
rect 20956 8792 24072 8820
rect 24171 8792 24216 8820
rect 20956 8780 20962 8792
rect 24210 8780 24216 8792
rect 24268 8780 24274 8832
rect 26602 8780 26608 8832
rect 26660 8820 26666 8832
rect 27433 8823 27491 8829
rect 27433 8820 27445 8823
rect 26660 8792 27445 8820
rect 26660 8780 26666 8792
rect 27433 8789 27445 8792
rect 27479 8789 27491 8823
rect 27433 8783 27491 8789
rect 1104 8730 38824 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 38824 8730
rect 1104 8656 38824 8678
rect 17310 8576 17316 8628
rect 17368 8616 17374 8628
rect 19165 8619 19223 8625
rect 19165 8616 19177 8619
rect 17368 8588 19177 8616
rect 17368 8576 17374 8588
rect 19165 8585 19177 8588
rect 19211 8585 19223 8619
rect 19165 8579 19223 8585
rect 20070 8576 20076 8628
rect 20128 8616 20134 8628
rect 21266 8616 21272 8628
rect 20128 8588 21272 8616
rect 20128 8576 20134 8588
rect 21266 8576 21272 8588
rect 21324 8616 21330 8628
rect 22186 8616 22192 8628
rect 21324 8588 22192 8616
rect 21324 8576 21330 8588
rect 22186 8576 22192 8588
rect 22244 8576 22250 8628
rect 22925 8619 22983 8625
rect 22925 8585 22937 8619
rect 22971 8616 22983 8619
rect 24854 8616 24860 8628
rect 22971 8588 24860 8616
rect 22971 8585 22983 8588
rect 22925 8579 22983 8585
rect 24854 8576 24860 8588
rect 24912 8576 24918 8628
rect 25774 8576 25780 8628
rect 25832 8616 25838 8628
rect 25869 8619 25927 8625
rect 25869 8616 25881 8619
rect 25832 8588 25881 8616
rect 25832 8576 25838 8588
rect 25869 8585 25881 8588
rect 25915 8585 25927 8619
rect 26510 8616 26516 8628
rect 26471 8588 26516 8616
rect 25869 8579 25927 8585
rect 26510 8576 26516 8588
rect 26568 8576 26574 8628
rect 27172 8588 27936 8616
rect 25590 8548 25596 8560
rect 24320 8520 25596 8548
rect 17954 8440 17960 8492
rect 18012 8480 18018 8492
rect 19889 8483 19947 8489
rect 19889 8480 19901 8483
rect 18012 8452 19901 8480
rect 18012 8440 18018 8452
rect 19889 8449 19901 8452
rect 19935 8449 19947 8483
rect 21637 8483 21695 8489
rect 21637 8480 21649 8483
rect 19889 8443 19947 8449
rect 19996 8452 21649 8480
rect 19426 8372 19432 8424
rect 19484 8412 19490 8424
rect 19996 8412 20024 8452
rect 21637 8449 21649 8452
rect 21683 8449 21695 8483
rect 21637 8443 21695 8449
rect 22922 8440 22928 8492
rect 22980 8480 22986 8492
rect 24320 8480 24348 8520
rect 25590 8508 25596 8520
rect 25648 8508 25654 8560
rect 22980 8452 24348 8480
rect 24765 8483 24823 8489
rect 22980 8440 22986 8452
rect 24765 8449 24777 8483
rect 24811 8480 24823 8483
rect 27172 8480 27200 8588
rect 24811 8452 27200 8480
rect 27908 8480 27936 8588
rect 28077 8483 28135 8489
rect 28077 8480 28089 8483
rect 27908 8452 28089 8480
rect 24811 8449 24823 8452
rect 24765 8443 24823 8449
rect 28077 8449 28089 8452
rect 28123 8449 28135 8483
rect 28077 8443 28135 8449
rect 19484 8384 20024 8412
rect 19484 8372 19490 8384
rect 22554 8372 22560 8424
rect 22612 8412 22618 8424
rect 23017 8415 23075 8421
rect 23017 8412 23029 8415
rect 22612 8384 23029 8412
rect 22612 8372 22618 8384
rect 23017 8381 23029 8384
rect 23063 8381 23075 8415
rect 25222 8412 25228 8424
rect 25183 8384 25228 8412
rect 23017 8375 23075 8381
rect 25222 8372 25228 8384
rect 25280 8372 25286 8424
rect 26053 8415 26111 8421
rect 26053 8412 26065 8415
rect 25424 8384 26065 8412
rect 18690 8304 18696 8356
rect 18748 8304 18754 8356
rect 20898 8304 20904 8356
rect 20956 8304 20962 8356
rect 21361 8347 21419 8353
rect 21361 8313 21373 8347
rect 21407 8344 21419 8347
rect 23293 8347 23351 8353
rect 21407 8316 23244 8344
rect 21407 8313 21419 8316
rect 21361 8307 21419 8313
rect 17678 8276 17684 8288
rect 17639 8248 17684 8276
rect 17678 8236 17684 8248
rect 17736 8236 17742 8288
rect 18782 8236 18788 8288
rect 18840 8276 18846 8288
rect 22925 8279 22983 8285
rect 22925 8276 22937 8279
rect 18840 8248 22937 8276
rect 18840 8236 18846 8248
rect 22925 8245 22937 8248
rect 22971 8245 22983 8279
rect 23216 8276 23244 8316
rect 23293 8313 23305 8347
rect 23339 8344 23351 8347
rect 23566 8344 23572 8356
rect 23339 8316 23572 8344
rect 23339 8313 23351 8316
rect 23293 8307 23351 8313
rect 23566 8304 23572 8316
rect 23624 8304 23630 8356
rect 25038 8344 25044 8356
rect 24518 8316 25044 8344
rect 25038 8304 25044 8316
rect 25096 8304 25102 8356
rect 25314 8276 25320 8288
rect 23216 8248 25320 8276
rect 22925 8239 22983 8245
rect 25314 8236 25320 8248
rect 25372 8236 25378 8288
rect 25424 8285 25452 8384
rect 26053 8381 26065 8384
rect 26099 8412 26111 8415
rect 26697 8415 26755 8421
rect 26697 8412 26709 8415
rect 26099 8384 26709 8412
rect 26099 8381 26111 8384
rect 26053 8375 26111 8381
rect 26697 8381 26709 8384
rect 26743 8412 26755 8415
rect 27338 8412 27344 8424
rect 26743 8384 27344 8412
rect 26743 8381 26755 8384
rect 26697 8375 26755 8381
rect 27338 8372 27344 8384
rect 27396 8372 27402 8424
rect 27801 8415 27859 8421
rect 27801 8381 27813 8415
rect 27847 8381 27859 8415
rect 27801 8375 27859 8381
rect 26786 8304 26792 8356
rect 26844 8344 26850 8356
rect 27816 8344 27844 8375
rect 29178 8372 29184 8424
rect 29236 8372 29242 8424
rect 30193 8415 30251 8421
rect 30193 8381 30205 8415
rect 30239 8412 30251 8415
rect 30374 8412 30380 8424
rect 30239 8384 30380 8412
rect 30239 8381 30251 8384
rect 30193 8375 30251 8381
rect 30374 8372 30380 8384
rect 30432 8412 30438 8424
rect 31478 8412 31484 8424
rect 30432 8384 31484 8412
rect 30432 8372 30438 8384
rect 31478 8372 31484 8384
rect 31536 8372 31542 8424
rect 26844 8316 27844 8344
rect 29380 8316 30052 8344
rect 26844 8304 26850 8316
rect 25409 8279 25467 8285
rect 25409 8245 25421 8279
rect 25455 8245 25467 8279
rect 25409 8239 25467 8245
rect 25774 8236 25780 8288
rect 25832 8276 25838 8288
rect 29380 8276 29408 8316
rect 29546 8276 29552 8288
rect 25832 8248 29408 8276
rect 29507 8248 29552 8276
rect 25832 8236 25838 8248
rect 29546 8236 29552 8248
rect 29604 8236 29610 8288
rect 30024 8285 30052 8316
rect 30009 8279 30067 8285
rect 30009 8245 30021 8279
rect 30055 8245 30067 8279
rect 30009 8239 30067 8245
rect 1104 8186 38824 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 38824 8186
rect 1104 8112 38824 8134
rect 19061 8075 19119 8081
rect 17328 8044 18920 8072
rect 16025 7939 16083 7945
rect 16025 7905 16037 7939
rect 16071 7905 16083 7939
rect 16025 7899 16083 7905
rect 14918 7760 14924 7812
rect 14976 7800 14982 7812
rect 16040 7800 16068 7899
rect 16206 7896 16212 7948
rect 16264 7936 16270 7948
rect 16853 7939 16911 7945
rect 16853 7936 16865 7939
rect 16264 7908 16865 7936
rect 16264 7896 16270 7908
rect 16853 7905 16865 7908
rect 16899 7936 16911 7939
rect 17218 7936 17224 7948
rect 16899 7908 17224 7936
rect 16899 7905 16911 7908
rect 16853 7899 16911 7905
rect 17218 7896 17224 7908
rect 17276 7896 17282 7948
rect 17328 7945 17356 8044
rect 17589 8007 17647 8013
rect 17589 7973 17601 8007
rect 17635 8004 17647 8007
rect 17678 8004 17684 8016
rect 17635 7976 17684 8004
rect 17635 7973 17647 7976
rect 17589 7967 17647 7973
rect 17678 7964 17684 7976
rect 17736 7964 17742 8016
rect 18892 8004 18920 8044
rect 19061 8041 19073 8075
rect 19107 8072 19119 8075
rect 20162 8072 20168 8084
rect 19107 8044 20168 8072
rect 19107 8041 19119 8044
rect 19061 8035 19119 8041
rect 20162 8032 20168 8044
rect 20220 8032 20226 8084
rect 20254 8032 20260 8084
rect 20312 8072 20318 8084
rect 23474 8072 23480 8084
rect 20312 8044 23480 8072
rect 20312 8032 20318 8044
rect 23474 8032 23480 8044
rect 23532 8032 23538 8084
rect 23566 8032 23572 8084
rect 23624 8072 23630 8084
rect 24305 8075 24363 8081
rect 24305 8072 24317 8075
rect 23624 8044 24317 8072
rect 23624 8032 23630 8044
rect 24305 8041 24317 8044
rect 24351 8041 24363 8075
rect 24305 8035 24363 8041
rect 26234 8032 26240 8084
rect 26292 8072 26298 8084
rect 27433 8075 27491 8081
rect 27433 8072 27445 8075
rect 26292 8044 27445 8072
rect 26292 8032 26298 8044
rect 27433 8041 27445 8044
rect 27479 8041 27491 8075
rect 30282 8072 30288 8084
rect 27433 8035 27491 8041
rect 27632 8044 30288 8072
rect 22922 8004 22928 8016
rect 18892 7976 19472 8004
rect 21850 7976 22928 8004
rect 19444 7948 19472 7976
rect 22922 7964 22928 7976
rect 22980 7964 22986 8016
rect 25774 8004 25780 8016
rect 24058 7976 25780 8004
rect 25774 7964 25780 7976
rect 25832 7964 25838 8016
rect 27632 8004 27660 8044
rect 30282 8032 30288 8044
rect 30340 8032 30346 8084
rect 31113 8075 31171 8081
rect 31113 8041 31125 8075
rect 31159 8041 31171 8075
rect 31113 8035 31171 8041
rect 26726 7976 27660 8004
rect 28905 8007 28963 8013
rect 28905 7973 28917 8007
rect 28951 8004 28963 8007
rect 29546 8004 29552 8016
rect 28951 7976 29552 8004
rect 28951 7973 28963 7976
rect 28905 7967 28963 7973
rect 29546 7964 29552 7976
rect 29604 7964 29610 8016
rect 31128 8004 31156 8035
rect 29656 7976 31156 8004
rect 17313 7939 17371 7945
rect 17313 7905 17325 7939
rect 17359 7905 17371 7939
rect 17313 7899 17371 7905
rect 18690 7896 18696 7948
rect 18748 7896 18754 7948
rect 19426 7896 19432 7948
rect 19484 7936 19490 7948
rect 19886 7936 19892 7948
rect 19484 7908 19892 7936
rect 19484 7896 19490 7908
rect 19886 7896 19892 7908
rect 19944 7936 19950 7948
rect 20349 7939 20407 7945
rect 20349 7936 20361 7939
rect 19944 7908 20361 7936
rect 19944 7896 19950 7908
rect 20349 7905 20361 7908
rect 20395 7905 20407 7939
rect 20349 7899 20407 7905
rect 27338 7896 27344 7948
rect 27396 7936 27402 7948
rect 29181 7939 29239 7945
rect 27396 7908 27830 7936
rect 27396 7896 27402 7908
rect 29181 7905 29193 7939
rect 29227 7936 29239 7939
rect 29270 7936 29276 7948
rect 29227 7908 29276 7936
rect 29227 7905 29239 7908
rect 29181 7899 29239 7905
rect 29270 7896 29276 7908
rect 29328 7936 29334 7948
rect 29656 7936 29684 7976
rect 29328 7908 29684 7936
rect 30653 7939 30711 7945
rect 29328 7896 29334 7908
rect 30653 7905 30665 7939
rect 30699 7905 30711 7939
rect 31294 7936 31300 7948
rect 31255 7908 31300 7936
rect 30653 7899 30711 7905
rect 19334 7868 19340 7880
rect 17420 7840 19340 7868
rect 17420 7800 17448 7840
rect 19334 7828 19340 7840
rect 19392 7828 19398 7880
rect 20625 7871 20683 7877
rect 20625 7837 20637 7871
rect 20671 7868 20683 7871
rect 22554 7868 22560 7880
rect 20671 7840 22094 7868
rect 22515 7840 22560 7868
rect 20671 7837 20683 7840
rect 20625 7831 20683 7837
rect 14976 7772 17448 7800
rect 22066 7800 22094 7840
rect 22554 7828 22560 7840
rect 22612 7828 22618 7880
rect 22830 7868 22836 7880
rect 22791 7840 22836 7868
rect 22830 7828 22836 7840
rect 22888 7828 22894 7880
rect 23474 7828 23480 7880
rect 23532 7868 23538 7880
rect 23532 7840 25084 7868
rect 23532 7828 23538 7840
rect 22066 7772 22692 7800
rect 14976 7760 14982 7772
rect 15102 7692 15108 7744
rect 15160 7732 15166 7744
rect 16209 7735 16267 7741
rect 16209 7732 16221 7735
rect 15160 7704 16221 7732
rect 15160 7692 15166 7704
rect 16209 7701 16221 7704
rect 16255 7701 16267 7735
rect 16666 7732 16672 7744
rect 16627 7704 16672 7732
rect 16209 7695 16267 7701
rect 16666 7692 16672 7704
rect 16724 7692 16730 7744
rect 16758 7692 16764 7744
rect 16816 7732 16822 7744
rect 20990 7732 20996 7744
rect 16816 7704 20996 7732
rect 16816 7692 16822 7704
rect 20990 7692 20996 7704
rect 21048 7692 21054 7744
rect 22097 7735 22155 7741
rect 22097 7701 22109 7735
rect 22143 7732 22155 7735
rect 22370 7732 22376 7744
rect 22143 7704 22376 7732
rect 22143 7701 22155 7704
rect 22097 7695 22155 7701
rect 22370 7692 22376 7704
rect 22428 7692 22434 7744
rect 22664 7732 22692 7772
rect 24946 7732 24952 7744
rect 22664 7704 24952 7732
rect 24946 7692 24952 7704
rect 25004 7692 25010 7744
rect 25056 7732 25084 7840
rect 25130 7828 25136 7880
rect 25188 7868 25194 7880
rect 25225 7871 25283 7877
rect 25225 7868 25237 7871
rect 25188 7840 25237 7868
rect 25188 7828 25194 7840
rect 25225 7837 25237 7840
rect 25271 7837 25283 7871
rect 25498 7868 25504 7880
rect 25459 7840 25504 7868
rect 25225 7831 25283 7837
rect 25498 7828 25504 7840
rect 25556 7828 25562 7880
rect 25590 7828 25596 7880
rect 25648 7868 25654 7880
rect 26973 7871 27031 7877
rect 26973 7868 26985 7871
rect 25648 7840 26985 7868
rect 25648 7828 25654 7840
rect 26973 7837 26985 7840
rect 27019 7837 27031 7871
rect 26973 7831 27031 7837
rect 28902 7828 28908 7880
rect 28960 7868 28966 7880
rect 28960 7840 29132 7868
rect 28960 7828 28966 7840
rect 29104 7800 29132 7840
rect 30668 7800 30696 7899
rect 31294 7896 31300 7908
rect 31352 7896 31358 7948
rect 29104 7772 30696 7800
rect 26602 7732 26608 7744
rect 25056 7704 26608 7732
rect 26602 7692 26608 7704
rect 26660 7692 26666 7744
rect 26786 7692 26792 7744
rect 26844 7732 26850 7744
rect 30469 7735 30527 7741
rect 30469 7732 30481 7735
rect 26844 7704 30481 7732
rect 26844 7692 26850 7704
rect 30469 7701 30481 7704
rect 30515 7701 30527 7735
rect 30469 7695 30527 7701
rect 1104 7642 38824 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 38824 7642
rect 1104 7568 38824 7590
rect 16393 7531 16451 7537
rect 16393 7497 16405 7531
rect 16439 7528 16451 7531
rect 16758 7528 16764 7540
rect 16439 7500 16764 7528
rect 16439 7497 16451 7500
rect 16393 7491 16451 7497
rect 16758 7488 16764 7500
rect 16816 7488 16822 7540
rect 22741 7531 22799 7537
rect 19306 7500 21220 7528
rect 15105 7463 15163 7469
rect 15105 7429 15117 7463
rect 15151 7460 15163 7463
rect 16574 7460 16580 7472
rect 15151 7432 16580 7460
rect 15151 7429 15163 7432
rect 15105 7423 15163 7429
rect 16574 7420 16580 7432
rect 16632 7460 16638 7472
rect 16632 7432 17724 7460
rect 16632 7420 16638 7432
rect 15194 7352 15200 7404
rect 15252 7392 15258 7404
rect 17696 7401 17724 7432
rect 17681 7395 17739 7401
rect 15252 7364 16252 7392
rect 15252 7352 15258 7364
rect 16224 7336 16252 7364
rect 17681 7361 17693 7395
rect 17727 7361 17739 7395
rect 17681 7355 17739 7361
rect 17957 7395 18015 7401
rect 17957 7361 17969 7395
rect 18003 7392 18015 7395
rect 19306 7392 19334 7500
rect 21192 7460 21220 7500
rect 22741 7497 22753 7531
rect 22787 7528 22799 7531
rect 22830 7528 22836 7540
rect 22787 7500 22836 7528
rect 22787 7497 22799 7500
rect 22741 7491 22799 7497
rect 22830 7488 22836 7500
rect 22888 7488 22894 7540
rect 24118 7528 24124 7540
rect 22940 7500 24124 7528
rect 22940 7460 22968 7500
rect 24118 7488 24124 7500
rect 24176 7488 24182 7540
rect 24946 7528 24952 7540
rect 24907 7500 24952 7528
rect 24946 7488 24952 7500
rect 25004 7488 25010 7540
rect 25314 7488 25320 7540
rect 25372 7528 25378 7540
rect 28626 7528 28632 7540
rect 25372 7500 28632 7528
rect 25372 7488 25378 7500
rect 28626 7488 28632 7500
rect 28684 7488 28690 7540
rect 29178 7488 29184 7540
rect 29236 7528 29242 7540
rect 31297 7531 31355 7537
rect 31297 7528 31309 7531
rect 29236 7500 31309 7528
rect 29236 7488 29242 7500
rect 31297 7497 31309 7500
rect 31343 7497 31355 7531
rect 31297 7491 31355 7497
rect 30190 7460 30196 7472
rect 21192 7432 22968 7460
rect 30151 7432 30196 7460
rect 30190 7420 30196 7432
rect 30248 7420 30254 7472
rect 18003 7364 19334 7392
rect 18003 7361 18015 7364
rect 17957 7355 18015 7361
rect 19426 7352 19432 7404
rect 19484 7392 19490 7404
rect 20165 7395 20223 7401
rect 20165 7392 20177 7395
rect 19484 7364 20177 7392
rect 19484 7352 19490 7364
rect 20165 7361 20177 7364
rect 20211 7361 20223 7395
rect 20165 7355 20223 7361
rect 20530 7352 20536 7404
rect 20588 7392 20594 7404
rect 23658 7392 23664 7404
rect 20588 7364 23664 7392
rect 20588 7352 20594 7364
rect 23658 7352 23664 7364
rect 23716 7352 23722 7404
rect 24210 7392 24216 7404
rect 24171 7364 24216 7392
rect 24210 7352 24216 7364
rect 24268 7352 24274 7404
rect 24486 7392 24492 7404
rect 24447 7364 24492 7392
rect 24486 7352 24492 7364
rect 24544 7352 24550 7404
rect 25406 7352 25412 7404
rect 25464 7392 25470 7404
rect 26421 7395 26479 7401
rect 26421 7392 26433 7395
rect 25464 7364 26433 7392
rect 25464 7352 25470 7364
rect 26421 7361 26433 7364
rect 26467 7361 26479 7395
rect 26694 7392 26700 7404
rect 26655 7364 26700 7392
rect 26421 7355 26479 7361
rect 26694 7352 26700 7364
rect 26752 7352 26758 7404
rect 27706 7352 27712 7404
rect 27764 7392 27770 7404
rect 28077 7395 28135 7401
rect 28077 7392 28089 7395
rect 27764 7364 28089 7392
rect 27764 7352 27770 7364
rect 28077 7361 28089 7364
rect 28123 7361 28135 7395
rect 28077 7355 28135 7361
rect 28166 7352 28172 7404
rect 28224 7392 28230 7404
rect 29270 7392 29276 7404
rect 28224 7364 29276 7392
rect 28224 7352 28230 7364
rect 29270 7352 29276 7364
rect 29328 7392 29334 7404
rect 29546 7392 29552 7404
rect 29328 7364 29552 7392
rect 29328 7352 29334 7364
rect 29546 7352 29552 7364
rect 29604 7352 29610 7404
rect 14918 7324 14924 7336
rect 14879 7296 14924 7324
rect 14918 7284 14924 7296
rect 14976 7284 14982 7336
rect 15010 7284 15016 7336
rect 15068 7324 15074 7336
rect 15565 7327 15623 7333
rect 15565 7324 15577 7327
rect 15068 7296 15577 7324
rect 15068 7284 15074 7296
rect 15565 7293 15577 7296
rect 15611 7293 15623 7327
rect 16206 7324 16212 7336
rect 16167 7296 16212 7324
rect 15565 7287 15623 7293
rect 15580 7256 15608 7287
rect 16206 7284 16212 7296
rect 16264 7284 16270 7336
rect 19886 7324 19892 7336
rect 19847 7296 19892 7324
rect 19886 7284 19892 7296
rect 19944 7284 19950 7336
rect 26712 7324 26740 7352
rect 27801 7327 27859 7333
rect 27801 7324 27813 7327
rect 26712 7296 27813 7324
rect 27801 7293 27813 7296
rect 27847 7293 27859 7327
rect 30006 7324 30012 7336
rect 29967 7296 30012 7324
rect 27801 7287 27859 7293
rect 17862 7256 17868 7268
rect 15580 7228 17868 7256
rect 17862 7216 17868 7228
rect 17920 7216 17926 7268
rect 20438 7256 20444 7268
rect 19182 7228 20444 7256
rect 20438 7216 20444 7228
rect 20496 7216 20502 7268
rect 22646 7256 22652 7268
rect 21390 7228 22652 7256
rect 22646 7216 22652 7228
rect 22704 7216 22710 7268
rect 23782 7228 25176 7256
rect 15749 7191 15807 7197
rect 15749 7157 15761 7191
rect 15795 7188 15807 7191
rect 17494 7188 17500 7200
rect 15795 7160 17500 7188
rect 15795 7157 15807 7160
rect 15749 7151 15807 7157
rect 17494 7148 17500 7160
rect 17552 7148 17558 7200
rect 19429 7191 19487 7197
rect 19429 7157 19441 7191
rect 19475 7188 19487 7191
rect 19978 7188 19984 7200
rect 19475 7160 19984 7188
rect 19475 7157 19487 7160
rect 19429 7151 19487 7157
rect 19978 7148 19984 7160
rect 20036 7148 20042 7200
rect 21634 7188 21640 7200
rect 21595 7160 21640 7188
rect 21634 7148 21640 7160
rect 21692 7148 21698 7200
rect 25148 7188 25176 7228
rect 25958 7216 25964 7268
rect 26016 7216 26022 7268
rect 27816 7256 27844 7287
rect 30006 7284 30012 7296
rect 30064 7284 30070 7336
rect 30834 7324 30840 7336
rect 30795 7296 30840 7324
rect 30834 7284 30840 7296
rect 30892 7284 30898 7336
rect 31478 7324 31484 7336
rect 31439 7296 31484 7324
rect 31478 7284 31484 7296
rect 31536 7284 31542 7336
rect 28166 7256 28172 7268
rect 27816 7228 28172 7256
rect 28166 7216 28172 7228
rect 28224 7216 28230 7268
rect 29822 7256 29828 7268
rect 29302 7228 29828 7256
rect 29822 7216 29828 7228
rect 29880 7216 29886 7268
rect 27154 7188 27160 7200
rect 25148 7160 27160 7188
rect 27154 7148 27160 7160
rect 27212 7148 27218 7200
rect 28718 7148 28724 7200
rect 28776 7188 28782 7200
rect 29549 7191 29607 7197
rect 29549 7188 29561 7191
rect 28776 7160 29561 7188
rect 28776 7148 28782 7160
rect 29549 7157 29561 7160
rect 29595 7157 29607 7191
rect 29549 7151 29607 7157
rect 30374 7148 30380 7200
rect 30432 7188 30438 7200
rect 30653 7191 30711 7197
rect 30653 7188 30665 7191
rect 30432 7160 30665 7188
rect 30432 7148 30438 7160
rect 30653 7157 30665 7160
rect 30699 7157 30711 7191
rect 30653 7151 30711 7157
rect 1104 7098 38824 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 38824 7098
rect 1104 7024 38824 7046
rect 15102 6944 15108 6996
rect 15160 6984 15166 6996
rect 20162 6984 20168 6996
rect 15160 6956 16712 6984
rect 20123 6956 20168 6984
rect 15160 6944 15166 6956
rect 16022 6876 16028 6928
rect 16080 6876 16086 6928
rect 14642 6808 14648 6860
rect 14700 6848 14706 6860
rect 15102 6848 15108 6860
rect 14700 6820 15108 6848
rect 14700 6808 14706 6820
rect 15102 6808 15108 6820
rect 15160 6808 15166 6860
rect 16684 6848 16712 6956
rect 20162 6944 20168 6956
rect 20220 6944 20226 6996
rect 21192 6956 23520 6984
rect 20254 6916 20260 6928
rect 18814 6888 20260 6916
rect 20254 6876 20260 6888
rect 20312 6876 20318 6928
rect 21192 6902 21220 6956
rect 21634 6916 21640 6928
rect 21595 6888 21640 6916
rect 21634 6876 21640 6888
rect 21692 6876 21698 6928
rect 23290 6876 23296 6928
rect 23348 6876 23354 6928
rect 23492 6916 23520 6956
rect 24118 6944 24124 6996
rect 24176 6984 24182 6996
rect 29181 6987 29239 6993
rect 29181 6984 29193 6987
rect 24176 6956 29193 6984
rect 24176 6944 24182 6956
rect 29181 6953 29193 6956
rect 29227 6953 29239 6987
rect 30469 6987 30527 6993
rect 30469 6984 30481 6987
rect 29181 6947 29239 6953
rect 29288 6956 30481 6984
rect 25314 6916 25320 6928
rect 23492 6888 25320 6916
rect 25314 6876 25320 6888
rect 25372 6876 25378 6928
rect 25682 6876 25688 6928
rect 25740 6876 25746 6928
rect 26694 6876 26700 6928
rect 26752 6916 26758 6928
rect 27709 6919 27767 6925
rect 26752 6888 27016 6916
rect 26752 6876 26758 6888
rect 16758 6848 16764 6860
rect 16684 6820 16764 6848
rect 16758 6808 16764 6820
rect 16816 6808 16822 6860
rect 21913 6851 21971 6857
rect 21913 6817 21925 6851
rect 21959 6848 21971 6851
rect 22554 6848 22560 6860
rect 21959 6820 22560 6848
rect 21959 6817 21971 6820
rect 21913 6811 21971 6817
rect 22554 6808 22560 6820
rect 22612 6808 22618 6860
rect 24121 6851 24179 6857
rect 24121 6817 24133 6851
rect 24167 6848 24179 6851
rect 24394 6848 24400 6860
rect 24167 6820 24400 6848
rect 24167 6817 24179 6820
rect 24121 6811 24179 6817
rect 24394 6808 24400 6820
rect 24452 6808 24458 6860
rect 26988 6857 27016 6888
rect 27709 6885 27721 6919
rect 27755 6916 27767 6919
rect 27798 6916 27804 6928
rect 27755 6888 27804 6916
rect 27755 6885 27767 6888
rect 27709 6879 27767 6885
rect 27798 6876 27804 6888
rect 27856 6876 27862 6928
rect 29288 6916 29316 6956
rect 30469 6953 30481 6956
rect 30515 6953 30527 6987
rect 30469 6947 30527 6953
rect 28934 6888 29316 6916
rect 30006 6876 30012 6928
rect 30064 6916 30070 6928
rect 30064 6888 30788 6916
rect 30064 6876 30070 6888
rect 26973 6851 27031 6857
rect 26973 6817 26985 6851
rect 27019 6848 27031 6851
rect 27430 6848 27436 6860
rect 27019 6820 27436 6848
rect 27019 6817 27031 6820
rect 26973 6811 27031 6817
rect 27430 6808 27436 6820
rect 27488 6808 27494 6860
rect 30466 6808 30472 6860
rect 30524 6848 30530 6860
rect 30653 6851 30711 6857
rect 30653 6848 30665 6851
rect 30524 6820 30665 6848
rect 30524 6808 30530 6820
rect 30653 6817 30665 6820
rect 30699 6817 30711 6851
rect 30760 6848 30788 6888
rect 31294 6876 31300 6928
rect 31352 6916 31358 6928
rect 31352 6888 32076 6916
rect 31352 6876 31358 6888
rect 31113 6851 31171 6857
rect 31113 6848 31125 6851
rect 30760 6820 31125 6848
rect 30653 6811 30711 6817
rect 31113 6817 31125 6820
rect 31159 6817 31171 6851
rect 31113 6811 31171 6817
rect 31941 6851 31999 6857
rect 31941 6817 31953 6851
rect 31987 6817 31999 6851
rect 32048 6848 32076 6888
rect 32585 6851 32643 6857
rect 32585 6848 32597 6851
rect 32048 6820 32597 6848
rect 31941 6811 31999 6817
rect 32585 6817 32597 6820
rect 32631 6817 32643 6851
rect 32585 6811 32643 6817
rect 15378 6780 15384 6792
rect 15339 6752 15384 6780
rect 15378 6740 15384 6752
rect 15436 6740 15442 6792
rect 16574 6740 16580 6792
rect 16632 6780 16638 6792
rect 17313 6783 17371 6789
rect 17313 6780 17325 6783
rect 16632 6752 17325 6780
rect 16632 6740 16638 6752
rect 17313 6749 17325 6752
rect 17359 6749 17371 6783
rect 17313 6743 17371 6749
rect 17589 6783 17647 6789
rect 17589 6749 17601 6783
rect 17635 6780 17647 6783
rect 19061 6783 19119 6789
rect 17635 6752 19012 6780
rect 17635 6749 17647 6752
rect 17589 6743 17647 6749
rect 18984 6712 19012 6752
rect 19061 6749 19073 6783
rect 19107 6780 19119 6783
rect 22462 6780 22468 6792
rect 19107 6752 22468 6780
rect 19107 6749 19119 6752
rect 19061 6743 19119 6749
rect 22462 6740 22468 6752
rect 22520 6740 22526 6792
rect 23842 6780 23848 6792
rect 23803 6752 23848 6780
rect 23842 6740 23848 6752
rect 23900 6740 23906 6792
rect 24946 6740 24952 6792
rect 25004 6780 25010 6792
rect 26697 6783 26755 6789
rect 26697 6780 26709 6783
rect 25004 6752 26709 6780
rect 25004 6740 25010 6752
rect 26697 6749 26709 6752
rect 26743 6749 26755 6783
rect 31956 6780 31984 6811
rect 26697 6743 26755 6749
rect 27540 6752 31984 6780
rect 20622 6712 20628 6724
rect 18984 6684 20628 6712
rect 20622 6672 20628 6684
rect 20680 6672 20686 6724
rect 22373 6715 22431 6721
rect 22373 6681 22385 6715
rect 22419 6712 22431 6715
rect 22738 6712 22744 6724
rect 22419 6684 22744 6712
rect 22419 6681 22431 6684
rect 22373 6675 22431 6681
rect 22738 6672 22744 6684
rect 22796 6672 22802 6724
rect 27246 6672 27252 6724
rect 27304 6712 27310 6724
rect 27540 6712 27568 6752
rect 31757 6715 31815 6721
rect 31757 6712 31769 6715
rect 27304 6684 27568 6712
rect 28736 6684 30420 6712
rect 27304 6672 27310 6684
rect 16850 6644 16856 6656
rect 16811 6616 16856 6644
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 16942 6604 16948 6656
rect 17000 6644 17006 6656
rect 21174 6644 21180 6656
rect 17000 6616 21180 6644
rect 17000 6604 17006 6616
rect 21174 6604 21180 6616
rect 21232 6604 21238 6656
rect 22830 6604 22836 6656
rect 22888 6644 22894 6656
rect 25225 6647 25283 6653
rect 25225 6644 25237 6647
rect 22888 6616 25237 6644
rect 22888 6604 22894 6616
rect 25225 6613 25237 6616
rect 25271 6613 25283 6647
rect 25225 6607 25283 6613
rect 26142 6604 26148 6656
rect 26200 6644 26206 6656
rect 28736 6644 28764 6684
rect 26200 6616 28764 6644
rect 26200 6604 26206 6616
rect 28810 6604 28816 6656
rect 28868 6644 28874 6656
rect 29362 6644 29368 6656
rect 28868 6616 29368 6644
rect 28868 6604 28874 6616
rect 29362 6604 29368 6616
rect 29420 6604 29426 6656
rect 30392 6644 30420 6684
rect 30576 6684 31769 6712
rect 30576 6644 30604 6684
rect 31757 6681 31769 6684
rect 31803 6681 31815 6715
rect 31757 6675 31815 6681
rect 30392 6616 30604 6644
rect 30834 6604 30840 6656
rect 30892 6644 30898 6656
rect 31297 6647 31355 6653
rect 31297 6644 31309 6647
rect 30892 6616 31309 6644
rect 30892 6604 30898 6616
rect 31297 6613 31309 6616
rect 31343 6644 31355 6647
rect 31662 6644 31668 6656
rect 31343 6616 31668 6644
rect 31343 6613 31355 6616
rect 31297 6607 31355 6613
rect 31662 6604 31668 6616
rect 31720 6604 31726 6656
rect 32398 6644 32404 6656
rect 32359 6616 32404 6644
rect 32398 6604 32404 6616
rect 32456 6604 32462 6656
rect 1104 6554 38824 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 38824 6554
rect 1104 6480 38824 6502
rect 14645 6443 14703 6449
rect 14645 6409 14657 6443
rect 14691 6440 14703 6443
rect 15378 6440 15384 6452
rect 14691 6412 15384 6440
rect 14691 6409 14703 6412
rect 14645 6403 14703 6409
rect 15378 6400 15384 6412
rect 15436 6400 15442 6452
rect 16850 6400 16856 6452
rect 16908 6440 16914 6452
rect 16908 6412 22094 6440
rect 16908 6400 16914 6412
rect 14185 6375 14243 6381
rect 14185 6341 14197 6375
rect 14231 6341 14243 6375
rect 16942 6372 16948 6384
rect 14185 6335 14243 6341
rect 16316 6344 16948 6372
rect 14200 6304 14228 6335
rect 16022 6304 16028 6316
rect 14200 6276 16028 6304
rect 16022 6264 16028 6276
rect 16080 6264 16086 6316
rect 16117 6307 16175 6313
rect 16117 6273 16129 6307
rect 16163 6304 16175 6307
rect 16316 6304 16344 6344
rect 16942 6332 16948 6344
rect 17000 6332 17006 6384
rect 19426 6372 19432 6384
rect 19387 6344 19432 6372
rect 19426 6332 19432 6344
rect 19484 6332 19490 6384
rect 22066 6372 22094 6412
rect 22186 6400 22192 6452
rect 22244 6440 22250 6452
rect 24302 6440 24308 6452
rect 22244 6412 23888 6440
rect 24263 6412 24308 6440
rect 22244 6400 22250 6412
rect 22066 6344 22324 6372
rect 16163 6276 16344 6304
rect 16393 6307 16451 6313
rect 16163 6273 16175 6276
rect 16117 6267 16175 6273
rect 16393 6273 16405 6307
rect 16439 6304 16451 6307
rect 16574 6304 16580 6316
rect 16439 6276 16580 6304
rect 16439 6273 16451 6276
rect 16393 6267 16451 6273
rect 16574 6264 16580 6276
rect 16632 6304 16638 6316
rect 17681 6307 17739 6313
rect 17681 6304 17693 6307
rect 16632 6276 17693 6304
rect 16632 6264 16638 6276
rect 17681 6273 17693 6276
rect 17727 6273 17739 6307
rect 17954 6304 17960 6316
rect 17915 6276 17960 6304
rect 17681 6267 17739 6273
rect 14001 6239 14059 6245
rect 14001 6205 14013 6239
rect 14047 6205 14059 6239
rect 14001 6199 14059 6205
rect 14016 6100 14044 6199
rect 15194 6100 15200 6112
rect 14016 6072 15200 6100
rect 15194 6060 15200 6072
rect 15252 6060 15258 6112
rect 15672 6100 15700 6154
rect 16666 6100 16672 6112
rect 15672 6072 16672 6100
rect 16666 6060 16672 6072
rect 16724 6060 16730 6112
rect 17696 6100 17724 6267
rect 17954 6264 17960 6276
rect 18012 6264 18018 6316
rect 19150 6264 19156 6316
rect 19208 6304 19214 6316
rect 21637 6307 21695 6313
rect 21637 6304 21649 6307
rect 19208 6276 21649 6304
rect 19208 6264 19214 6276
rect 21637 6273 21649 6276
rect 21683 6273 21695 6307
rect 21637 6267 21695 6273
rect 19886 6236 19892 6248
rect 19847 6208 19892 6236
rect 19886 6196 19892 6208
rect 19944 6196 19950 6248
rect 21450 6196 21456 6248
rect 21508 6236 21514 6248
rect 22186 6236 22192 6248
rect 21508 6208 22192 6236
rect 21508 6196 21514 6208
rect 22186 6196 22192 6208
rect 22244 6196 22250 6248
rect 22296 6236 22324 6344
rect 22370 6264 22376 6316
rect 22428 6304 22434 6316
rect 22833 6307 22891 6313
rect 22833 6304 22845 6307
rect 22428 6276 22845 6304
rect 22428 6264 22434 6276
rect 22833 6273 22845 6276
rect 22879 6273 22891 6307
rect 23860 6304 23888 6412
rect 24302 6400 24308 6412
rect 24360 6400 24366 6452
rect 24854 6400 24860 6452
rect 24912 6440 24918 6452
rect 26786 6440 26792 6452
rect 24912 6412 26792 6440
rect 24912 6400 24918 6412
rect 26786 6400 26792 6412
rect 26844 6400 26850 6452
rect 27246 6400 27252 6452
rect 27304 6440 27310 6452
rect 27304 6412 29132 6440
rect 27304 6400 27310 6412
rect 29104 6372 29132 6412
rect 29822 6400 29828 6452
rect 29880 6440 29886 6452
rect 30009 6443 30067 6449
rect 30009 6440 30021 6443
rect 29880 6412 30021 6440
rect 29880 6400 29886 6412
rect 30009 6409 30021 6412
rect 30055 6409 30067 6443
rect 30009 6403 30067 6409
rect 30282 6400 30288 6452
rect 30340 6440 30346 6452
rect 31297 6443 31355 6449
rect 31297 6440 31309 6443
rect 30340 6412 31309 6440
rect 30340 6400 30346 6412
rect 31297 6409 31309 6412
rect 31343 6409 31355 6443
rect 31297 6403 31355 6409
rect 30466 6372 30472 6384
rect 29104 6344 30472 6372
rect 30466 6332 30472 6344
rect 30524 6332 30530 6384
rect 23860 6276 30880 6304
rect 22833 6267 22891 6273
rect 22554 6236 22560 6248
rect 22296 6208 22416 6236
rect 22515 6208 22560 6236
rect 19182 6140 20116 6168
rect 19334 6100 19340 6112
rect 17696 6072 19340 6100
rect 19334 6060 19340 6072
rect 19392 6060 19398 6112
rect 20088 6100 20116 6140
rect 20162 6128 20168 6180
rect 20220 6168 20226 6180
rect 20220 6140 20265 6168
rect 21390 6140 21588 6168
rect 20220 6128 20226 6140
rect 21450 6100 21456 6112
rect 20088 6072 21456 6100
rect 21450 6060 21456 6072
rect 21508 6060 21514 6112
rect 21560 6100 21588 6140
rect 21818 6128 21824 6180
rect 21876 6168 21882 6180
rect 22278 6168 22284 6180
rect 21876 6140 22284 6168
rect 21876 6128 21882 6140
rect 22278 6128 22284 6140
rect 22336 6128 22342 6180
rect 22094 6100 22100 6112
rect 21560 6072 22100 6100
rect 22094 6060 22100 6072
rect 22152 6060 22158 6112
rect 22388 6100 22416 6208
rect 22554 6196 22560 6208
rect 22612 6196 22618 6248
rect 24854 6236 24860 6248
rect 23966 6208 24860 6236
rect 24854 6196 24860 6208
rect 24912 6196 24918 6248
rect 26510 6196 26516 6248
rect 26568 6236 26574 6248
rect 26568 6208 26613 6236
rect 26568 6196 26574 6208
rect 27430 6196 27436 6248
rect 27488 6236 27494 6248
rect 27801 6239 27859 6245
rect 27801 6236 27813 6239
rect 27488 6208 27813 6236
rect 27488 6196 27494 6208
rect 27801 6205 27813 6208
rect 27847 6205 27859 6239
rect 27801 6199 27859 6205
rect 29362 6196 29368 6248
rect 29420 6236 29426 6248
rect 30193 6239 30251 6245
rect 30193 6236 30205 6239
rect 29420 6208 30205 6236
rect 29420 6196 29426 6208
rect 30193 6205 30205 6208
rect 30239 6205 30251 6239
rect 30193 6199 30251 6205
rect 30282 6196 30288 6248
rect 30340 6236 30346 6248
rect 30852 6245 30880 6276
rect 30837 6239 30895 6245
rect 30340 6208 30788 6236
rect 30340 6196 30346 6208
rect 26142 6168 26148 6180
rect 24136 6140 24900 6168
rect 25806 6140 26148 6168
rect 24136 6100 24164 6140
rect 24762 6100 24768 6112
rect 22388 6072 24164 6100
rect 24723 6072 24768 6100
rect 24762 6060 24768 6072
rect 24820 6060 24826 6112
rect 24872 6100 24900 6140
rect 26142 6128 26148 6140
rect 26200 6128 26206 6180
rect 26237 6171 26295 6177
rect 26237 6137 26249 6171
rect 26283 6168 26295 6171
rect 26970 6168 26976 6180
rect 26283 6140 26976 6168
rect 26283 6137 26295 6140
rect 26237 6131 26295 6137
rect 26970 6128 26976 6140
rect 27028 6128 27034 6180
rect 28077 6171 28135 6177
rect 28077 6137 28089 6171
rect 28123 6137 28135 6171
rect 30760 6168 30788 6208
rect 30837 6205 30849 6239
rect 30883 6205 30895 6239
rect 30837 6199 30895 6205
rect 31481 6239 31539 6245
rect 31481 6205 31493 6239
rect 31527 6205 31539 6239
rect 31481 6199 31539 6205
rect 32125 6239 32183 6245
rect 32125 6205 32137 6239
rect 32171 6205 32183 6239
rect 32125 6199 32183 6205
rect 31496 6168 31524 6199
rect 29302 6140 30696 6168
rect 30760 6140 31524 6168
rect 28077 6131 28135 6137
rect 28092 6100 28120 6131
rect 24872 6072 28120 6100
rect 28166 6060 28172 6112
rect 28224 6100 28230 6112
rect 30668 6109 30696 6140
rect 31662 6128 31668 6180
rect 31720 6168 31726 6180
rect 32140 6168 32168 6199
rect 31720 6140 32168 6168
rect 31720 6128 31726 6140
rect 29549 6103 29607 6109
rect 29549 6100 29561 6103
rect 28224 6072 29561 6100
rect 28224 6060 28230 6072
rect 29549 6069 29561 6072
rect 29595 6069 29607 6103
rect 29549 6063 29607 6069
rect 30653 6103 30711 6109
rect 30653 6069 30665 6103
rect 30699 6069 30711 6103
rect 31938 6100 31944 6112
rect 31899 6072 31944 6100
rect 30653 6063 30711 6069
rect 31938 6060 31944 6072
rect 31996 6060 32002 6112
rect 1104 6010 38824 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 38824 6010
rect 1104 5936 38824 5958
rect 13817 5899 13875 5905
rect 13817 5865 13829 5899
rect 13863 5865 13875 5899
rect 17310 5896 17316 5908
rect 17271 5868 17316 5896
rect 13817 5859 13875 5865
rect 13832 5828 13860 5859
rect 17310 5856 17316 5868
rect 17368 5856 17374 5908
rect 21542 5896 21548 5908
rect 18340 5868 21548 5896
rect 13832 5800 15410 5828
rect 18340 5814 18368 5868
rect 21542 5856 21548 5868
rect 21600 5856 21606 5908
rect 24118 5896 24124 5908
rect 21744 5868 24124 5896
rect 21744 5814 21772 5868
rect 24118 5856 24124 5868
rect 24176 5856 24182 5908
rect 24213 5899 24271 5905
rect 24213 5865 24225 5899
rect 24259 5896 24271 5899
rect 25406 5896 25412 5908
rect 24259 5868 25412 5896
rect 24259 5865 24271 5868
rect 24213 5859 24271 5865
rect 25406 5856 25412 5868
rect 25464 5856 25470 5908
rect 26970 5896 26976 5908
rect 26931 5868 26976 5896
rect 26970 5856 26976 5868
rect 27028 5856 27034 5908
rect 30374 5896 30380 5908
rect 27632 5868 30380 5896
rect 22741 5831 22799 5837
rect 22741 5797 22753 5831
rect 22787 5828 22799 5831
rect 22830 5828 22836 5840
rect 22787 5800 22836 5828
rect 22787 5797 22799 5800
rect 22741 5791 22799 5797
rect 22830 5788 22836 5800
rect 22888 5788 22894 5840
rect 23750 5788 23756 5840
rect 23808 5788 23814 5840
rect 24854 5788 24860 5840
rect 24912 5828 24918 5840
rect 25501 5831 25559 5837
rect 25501 5828 25513 5831
rect 24912 5800 25513 5828
rect 24912 5788 24918 5800
rect 25501 5797 25513 5800
rect 25547 5797 25559 5831
rect 27632 5828 27660 5868
rect 30374 5856 30380 5868
rect 30432 5856 30438 5908
rect 26726 5800 27660 5828
rect 25501 5791 25559 5797
rect 28442 5788 28448 5840
rect 28500 5788 28506 5840
rect 28810 5788 28816 5840
rect 28868 5828 28874 5840
rect 28868 5800 31248 5828
rect 28868 5788 28874 5800
rect 13633 5763 13691 5769
rect 13633 5729 13645 5763
rect 13679 5760 13691 5763
rect 15010 5760 15016 5772
rect 13679 5732 15016 5760
rect 13679 5729 13691 5732
rect 13633 5723 13691 5729
rect 15010 5720 15016 5732
rect 15068 5720 15074 5772
rect 16850 5720 16856 5772
rect 16908 5760 16914 5772
rect 19061 5763 19119 5769
rect 16908 5732 16953 5760
rect 16908 5720 16914 5732
rect 19061 5729 19073 5763
rect 19107 5760 19119 5763
rect 19334 5760 19340 5772
rect 19107 5732 19340 5760
rect 19107 5729 19119 5732
rect 19061 5723 19119 5729
rect 19334 5720 19340 5732
rect 19392 5760 19398 5772
rect 20257 5763 20315 5769
rect 20257 5760 20269 5763
rect 19392 5732 20269 5760
rect 19392 5720 19398 5732
rect 20257 5729 20269 5732
rect 20303 5729 20315 5763
rect 22462 5760 22468 5772
rect 22423 5732 22468 5760
rect 20257 5723 20315 5729
rect 22462 5720 22468 5732
rect 22520 5720 22526 5772
rect 24394 5720 24400 5772
rect 24452 5760 24458 5772
rect 25222 5760 25228 5772
rect 24452 5732 25228 5760
rect 24452 5720 24458 5732
rect 25222 5720 25228 5732
rect 25280 5720 25286 5772
rect 29196 5769 29224 5800
rect 29181 5763 29239 5769
rect 29181 5729 29193 5763
rect 29227 5729 29239 5763
rect 29181 5723 29239 5729
rect 29270 5720 29276 5772
rect 29328 5760 29334 5772
rect 30653 5763 30711 5769
rect 30653 5760 30665 5763
rect 29328 5732 30665 5760
rect 29328 5720 29334 5732
rect 30653 5729 30665 5732
rect 30699 5729 30711 5763
rect 30653 5723 30711 5729
rect 31113 5763 31171 5769
rect 31113 5729 31125 5763
rect 31159 5729 31171 5763
rect 31113 5723 31171 5729
rect 16577 5695 16635 5701
rect 16577 5661 16589 5695
rect 16623 5692 16635 5695
rect 18782 5692 18788 5704
rect 16623 5664 16804 5692
rect 18743 5664 18788 5692
rect 16623 5661 16635 5664
rect 16577 5655 16635 5661
rect 16776 5624 16804 5664
rect 18782 5652 18788 5664
rect 18840 5652 18846 5704
rect 20533 5695 20591 5701
rect 20533 5661 20545 5695
rect 20579 5692 20591 5695
rect 22278 5692 22284 5704
rect 20579 5664 22284 5692
rect 20579 5661 20591 5664
rect 20533 5655 20591 5661
rect 22278 5652 22284 5664
rect 22336 5652 22342 5704
rect 28166 5692 28172 5704
rect 22572 5664 28172 5692
rect 22572 5624 22600 5664
rect 28166 5652 28172 5664
rect 28224 5652 28230 5704
rect 28350 5652 28356 5704
rect 28408 5692 28414 5704
rect 28905 5695 28963 5701
rect 28905 5692 28917 5695
rect 28408 5664 28917 5692
rect 28408 5652 28414 5664
rect 28905 5661 28917 5664
rect 28951 5661 28963 5695
rect 28905 5655 28963 5661
rect 30006 5652 30012 5704
rect 30064 5692 30070 5704
rect 31128 5692 31156 5723
rect 30064 5664 31156 5692
rect 31220 5692 31248 5800
rect 31386 5788 31392 5840
rect 31444 5828 31450 5840
rect 31662 5828 31668 5840
rect 31444 5800 31668 5828
rect 31444 5788 31450 5800
rect 31662 5788 31668 5800
rect 31720 5828 31726 5840
rect 31720 5800 32628 5828
rect 31720 5788 31726 5800
rect 31294 5720 31300 5772
rect 31352 5760 31358 5772
rect 32600 5769 32628 5800
rect 31941 5763 31999 5769
rect 31941 5760 31953 5763
rect 31352 5732 31953 5760
rect 31352 5720 31358 5732
rect 31941 5729 31953 5732
rect 31987 5729 31999 5763
rect 31941 5723 31999 5729
rect 32585 5763 32643 5769
rect 32585 5729 32597 5763
rect 32631 5729 32643 5763
rect 32585 5723 32643 5729
rect 32398 5692 32404 5704
rect 31220 5664 32404 5692
rect 30064 5652 30070 5664
rect 32398 5652 32404 5664
rect 32456 5652 32462 5704
rect 16776 5596 17816 5624
rect 15102 5556 15108 5568
rect 15063 5528 15108 5556
rect 15102 5516 15108 5528
rect 15160 5516 15166 5568
rect 17788 5556 17816 5596
rect 21560 5596 22600 5624
rect 27264 5596 27936 5624
rect 21560 5556 21588 5596
rect 17788 5528 21588 5556
rect 22005 5559 22063 5565
rect 22005 5525 22017 5559
rect 22051 5556 22063 5559
rect 22830 5556 22836 5568
rect 22051 5528 22836 5556
rect 22051 5525 22063 5528
rect 22005 5519 22063 5525
rect 22830 5516 22836 5528
rect 22888 5516 22894 5568
rect 24118 5516 24124 5568
rect 24176 5556 24182 5568
rect 27264 5556 27292 5596
rect 27430 5556 27436 5568
rect 24176 5528 27292 5556
rect 27391 5528 27436 5556
rect 24176 5516 24182 5528
rect 27430 5516 27436 5528
rect 27488 5516 27494 5568
rect 27908 5556 27936 5596
rect 29362 5584 29368 5636
rect 29420 5624 29426 5636
rect 30282 5624 30288 5636
rect 29420 5596 30288 5624
rect 29420 5584 29426 5596
rect 30282 5584 30288 5596
rect 30340 5584 30346 5636
rect 30392 5596 32444 5624
rect 28166 5556 28172 5568
rect 27908 5528 28172 5556
rect 28166 5516 28172 5528
rect 28224 5516 28230 5568
rect 28258 5516 28264 5568
rect 28316 5556 28322 5568
rect 30392 5556 30420 5596
rect 28316 5528 30420 5556
rect 28316 5516 28322 5528
rect 30466 5516 30472 5568
rect 30524 5556 30530 5568
rect 31294 5556 31300 5568
rect 30524 5528 30569 5556
rect 31255 5528 31300 5556
rect 30524 5516 30530 5528
rect 31294 5516 31300 5528
rect 31352 5516 31358 5568
rect 31754 5556 31760 5568
rect 31715 5528 31760 5556
rect 31754 5516 31760 5528
rect 31812 5516 31818 5568
rect 32416 5565 32444 5596
rect 32401 5559 32459 5565
rect 32401 5525 32413 5559
rect 32447 5525 32459 5559
rect 32401 5519 32459 5525
rect 1104 5466 38824 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 38824 5466
rect 1104 5392 38824 5414
rect 17681 5355 17739 5361
rect 17681 5321 17693 5355
rect 17727 5352 17739 5355
rect 18782 5352 18788 5364
rect 17727 5324 18788 5352
rect 17727 5321 17739 5324
rect 17681 5315 17739 5321
rect 18782 5312 18788 5324
rect 18840 5312 18846 5364
rect 24854 5352 24860 5364
rect 24815 5324 24860 5352
rect 24854 5312 24860 5324
rect 24912 5312 24918 5364
rect 30653 5355 30711 5361
rect 30653 5352 30665 5355
rect 25148 5324 30665 5352
rect 24397 5287 24455 5293
rect 24397 5253 24409 5287
rect 24443 5284 24455 5287
rect 24946 5284 24952 5296
rect 24443 5256 24952 5284
rect 24443 5253 24455 5256
rect 24397 5247 24455 5253
rect 24946 5244 24952 5256
rect 25004 5244 25010 5296
rect 14093 5219 14151 5225
rect 14093 5185 14105 5219
rect 14139 5216 14151 5219
rect 16482 5216 16488 5228
rect 14139 5188 16488 5216
rect 14139 5185 14151 5188
rect 14093 5179 14151 5185
rect 16482 5176 16488 5188
rect 16540 5176 16546 5228
rect 19426 5216 19432 5228
rect 19387 5188 19432 5216
rect 19426 5176 19432 5188
rect 19484 5216 19490 5228
rect 19889 5219 19947 5225
rect 19889 5216 19901 5219
rect 19484 5188 19901 5216
rect 19484 5176 19490 5188
rect 19889 5185 19901 5188
rect 19935 5185 19947 5219
rect 19889 5179 19947 5185
rect 20165 5219 20223 5225
rect 20165 5185 20177 5219
rect 20211 5216 20223 5219
rect 21174 5216 21180 5228
rect 20211 5188 21180 5216
rect 20211 5185 20223 5188
rect 20165 5179 20223 5185
rect 21174 5176 21180 5188
rect 21232 5176 21238 5228
rect 22554 5176 22560 5228
rect 22612 5216 22618 5228
rect 22649 5219 22707 5225
rect 22649 5216 22661 5219
rect 22612 5188 22661 5216
rect 22612 5176 22618 5188
rect 22649 5185 22661 5188
rect 22695 5185 22707 5219
rect 22649 5179 22707 5185
rect 22925 5219 22983 5225
rect 22925 5185 22937 5219
rect 22971 5216 22983 5219
rect 24762 5216 24768 5228
rect 22971 5188 24768 5216
rect 22971 5185 22983 5188
rect 22925 5179 22983 5185
rect 24762 5176 24768 5188
rect 24820 5176 24826 5228
rect 14185 5151 14243 5157
rect 14185 5117 14197 5151
rect 14231 5117 14243 5151
rect 14642 5148 14648 5160
rect 14603 5120 14648 5148
rect 14185 5111 14243 5117
rect 14200 5012 14228 5111
rect 14642 5108 14648 5120
rect 14700 5108 14706 5160
rect 21298 5120 22600 5148
rect 14918 5080 14924 5092
rect 14879 5052 14924 5080
rect 14918 5040 14924 5052
rect 14976 5040 14982 5092
rect 17862 5080 17868 5092
rect 16146 5052 17868 5080
rect 17862 5040 17868 5052
rect 17920 5040 17926 5092
rect 19058 5080 19064 5092
rect 18722 5052 19064 5080
rect 19058 5040 19064 5052
rect 19116 5040 19122 5092
rect 19153 5083 19211 5089
rect 19153 5049 19165 5083
rect 19199 5080 19211 5083
rect 20070 5080 20076 5092
rect 19199 5052 20076 5080
rect 19199 5049 19211 5052
rect 19153 5043 19211 5049
rect 20070 5040 20076 5052
rect 20128 5040 20134 5092
rect 15102 5012 15108 5024
rect 14200 4984 15108 5012
rect 15102 4972 15108 4984
rect 15160 4972 15166 5024
rect 16393 5015 16451 5021
rect 16393 4981 16405 5015
rect 16439 5012 16451 5015
rect 17586 5012 17592 5024
rect 16439 4984 17592 5012
rect 16439 4981 16451 4984
rect 16393 4975 16451 4981
rect 17586 4972 17592 4984
rect 17644 4972 17650 5024
rect 21637 5015 21695 5021
rect 21637 4981 21649 5015
rect 21683 5012 21695 5015
rect 22370 5012 22376 5024
rect 21683 4984 22376 5012
rect 21683 4981 21695 4984
rect 21637 4975 21695 4981
rect 22370 4972 22376 4984
rect 22428 4972 22434 5024
rect 22572 5012 22600 5120
rect 24026 5108 24032 5160
rect 24084 5108 24090 5160
rect 25148 5148 25176 5324
rect 30653 5321 30665 5324
rect 30699 5321 30711 5355
rect 30653 5315 30711 5321
rect 28258 5284 28264 5296
rect 26528 5256 28264 5284
rect 25866 5176 25872 5228
rect 25924 5216 25930 5228
rect 26528 5216 26556 5256
rect 28258 5244 28264 5256
rect 28316 5244 28322 5296
rect 30374 5244 30380 5296
rect 30432 5284 30438 5296
rect 31297 5287 31355 5293
rect 31297 5284 31309 5287
rect 30432 5256 31309 5284
rect 30432 5244 30438 5256
rect 31297 5253 31309 5256
rect 31343 5253 31355 5287
rect 31297 5247 31355 5253
rect 25924 5188 26556 5216
rect 26605 5219 26663 5225
rect 25924 5176 25930 5188
rect 26605 5185 26617 5219
rect 26651 5216 26663 5219
rect 26694 5216 26700 5228
rect 26651 5188 26700 5216
rect 26651 5185 26663 5188
rect 26605 5179 26663 5185
rect 26694 5176 26700 5188
rect 26752 5176 26758 5228
rect 31938 5216 31944 5228
rect 27724 5188 31944 5216
rect 24228 5120 25176 5148
rect 24228 5012 24256 5120
rect 26326 5080 26332 5092
rect 22572 4984 24256 5012
rect 25884 5012 25912 5066
rect 26287 5052 26332 5080
rect 26326 5040 26332 5052
rect 26384 5040 26390 5092
rect 27724 5012 27752 5188
rect 31938 5176 31944 5188
rect 31996 5176 32002 5228
rect 29546 5108 29552 5160
rect 29604 5148 29610 5160
rect 29604 5120 29649 5148
rect 29604 5108 29610 5120
rect 30006 5108 30012 5160
rect 30064 5148 30070 5160
rect 30193 5151 30251 5157
rect 30193 5148 30205 5151
rect 30064 5120 30205 5148
rect 30064 5108 30070 5120
rect 30193 5117 30205 5120
rect 30239 5117 30251 5151
rect 30193 5111 30251 5117
rect 30650 5108 30656 5160
rect 30708 5148 30714 5160
rect 30837 5151 30895 5157
rect 30837 5148 30849 5151
rect 30708 5120 30849 5148
rect 30708 5108 30714 5120
rect 30837 5117 30849 5120
rect 30883 5148 30895 5151
rect 31294 5148 31300 5160
rect 30883 5120 31300 5148
rect 30883 5117 30895 5120
rect 30837 5111 30895 5117
rect 31294 5108 31300 5120
rect 31352 5148 31358 5160
rect 31481 5151 31539 5157
rect 31481 5148 31493 5151
rect 31352 5120 31493 5148
rect 31352 5108 31358 5120
rect 31481 5117 31493 5120
rect 31527 5117 31539 5151
rect 31481 5111 31539 5117
rect 27982 5040 27988 5092
rect 28040 5080 28046 5092
rect 29270 5080 29276 5092
rect 28040 5052 28106 5080
rect 29231 5052 29276 5080
rect 28040 5040 28046 5052
rect 29270 5040 29276 5052
rect 29328 5040 29334 5092
rect 25884 4984 27752 5012
rect 27801 5015 27859 5021
rect 27801 4981 27813 5015
rect 27847 5012 27859 5015
rect 27890 5012 27896 5024
rect 27847 4984 27896 5012
rect 27847 4981 27859 4984
rect 27801 4975 27859 4981
rect 27890 4972 27896 4984
rect 27948 4972 27954 5024
rect 28902 4972 28908 5024
rect 28960 5012 28966 5024
rect 30009 5015 30067 5021
rect 30009 5012 30021 5015
rect 28960 4984 30021 5012
rect 28960 4972 28966 4984
rect 30009 4981 30021 4984
rect 30055 4981 30067 5015
rect 30009 4975 30067 4981
rect 1104 4922 38824 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 38824 4922
rect 1104 4848 38824 4870
rect 14918 4768 14924 4820
rect 14976 4808 14982 4820
rect 15105 4811 15163 4817
rect 15105 4808 15117 4811
rect 14976 4780 15117 4808
rect 14976 4768 14982 4780
rect 15105 4777 15117 4780
rect 15151 4777 15163 4811
rect 15105 4771 15163 4777
rect 17862 4768 17868 4820
rect 17920 4808 17926 4820
rect 27893 4811 27951 4817
rect 17920 4780 27384 4808
rect 17920 4768 17926 4780
rect 16114 4700 16120 4752
rect 16172 4700 16178 4752
rect 18322 4700 18328 4752
rect 18380 4700 18386 4752
rect 22830 4740 22836 4752
rect 16850 4632 16856 4684
rect 16908 4672 16914 4684
rect 17310 4672 17316 4684
rect 16908 4644 17316 4672
rect 16908 4632 16914 4644
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 16574 4604 16580 4616
rect 16535 4576 16580 4604
rect 16574 4564 16580 4576
rect 16632 4564 16638 4616
rect 17678 4564 17684 4616
rect 17736 4604 17742 4616
rect 20456 4604 20484 4726
rect 22791 4712 22836 4740
rect 22830 4700 22836 4712
rect 22888 4700 22894 4752
rect 25866 4740 25872 4752
rect 24058 4712 25872 4740
rect 25866 4700 25872 4712
rect 25924 4700 25930 4752
rect 26234 4700 26240 4752
rect 26292 4700 26298 4752
rect 27356 4740 27384 4780
rect 27893 4777 27905 4811
rect 27939 4808 27951 4811
rect 29270 4808 29276 4820
rect 27939 4780 29276 4808
rect 27939 4777 27951 4780
rect 27893 4771 27951 4777
rect 29270 4768 29276 4780
rect 29328 4768 29334 4820
rect 28445 4743 28503 4749
rect 27356 4712 27936 4740
rect 22554 4672 22560 4684
rect 22066 4644 22560 4672
rect 17736 4576 20484 4604
rect 17736 4564 17742 4576
rect 20714 4564 20720 4616
rect 20772 4604 20778 4616
rect 21453 4607 21511 4613
rect 21453 4604 21465 4607
rect 20772 4576 21465 4604
rect 20772 4564 20778 4576
rect 21453 4573 21465 4576
rect 21499 4573 21511 4607
rect 21453 4567 21511 4573
rect 21821 4607 21879 4613
rect 21821 4573 21833 4607
rect 21867 4604 21879 4607
rect 22066 4604 22094 4644
rect 22554 4632 22560 4644
rect 22612 4632 22618 4684
rect 27065 4675 27123 4681
rect 27065 4641 27077 4675
rect 27111 4672 27123 4675
rect 27798 4672 27804 4684
rect 27111 4644 27804 4672
rect 27111 4641 27123 4644
rect 27065 4635 27123 4641
rect 27798 4632 27804 4644
rect 27856 4632 27862 4684
rect 21867 4576 22094 4604
rect 24305 4607 24363 4613
rect 21867 4573 21879 4576
rect 21821 4567 21879 4573
rect 24305 4573 24317 4607
rect 24351 4604 24363 4607
rect 26694 4604 26700 4616
rect 24351 4576 26700 4604
rect 24351 4573 24363 4576
rect 24305 4567 24363 4573
rect 19061 4539 19119 4545
rect 19061 4505 19073 4539
rect 19107 4536 19119 4539
rect 20622 4536 20628 4548
rect 19107 4508 20628 4536
rect 19107 4505 19119 4508
rect 19061 4499 19119 4505
rect 20622 4496 20628 4508
rect 20680 4496 20686 4548
rect 17576 4471 17634 4477
rect 17576 4437 17588 4471
rect 17622 4468 17634 4471
rect 19886 4468 19892 4480
rect 17622 4440 19892 4468
rect 17622 4437 17634 4440
rect 17576 4431 17634 4437
rect 19886 4428 19892 4440
rect 19944 4428 19950 4480
rect 19978 4428 19984 4480
rect 20036 4477 20042 4480
rect 20036 4471 20085 4477
rect 20036 4437 20039 4471
rect 20073 4437 20085 4471
rect 20036 4431 20085 4437
rect 20036 4428 20042 4431
rect 20438 4428 20444 4480
rect 20496 4468 20502 4480
rect 21836 4468 21864 4567
rect 26694 4564 26700 4576
rect 26752 4564 26758 4616
rect 26786 4564 26792 4616
rect 26844 4604 26850 4616
rect 27433 4607 27491 4613
rect 27433 4604 27445 4607
rect 26844 4576 27445 4604
rect 26844 4564 26850 4576
rect 27433 4573 27445 4576
rect 27479 4573 27491 4607
rect 27433 4567 27491 4573
rect 27908 4536 27936 4712
rect 28445 4709 28457 4743
rect 28491 4740 28503 4743
rect 28718 4740 28724 4752
rect 28491 4712 28724 4740
rect 28491 4709 28503 4712
rect 28445 4703 28503 4709
rect 28169 4675 28227 4681
rect 28169 4641 28181 4675
rect 28215 4672 28227 4675
rect 28460 4672 28488 4703
rect 28718 4700 28724 4712
rect 28776 4700 28782 4752
rect 29178 4672 29184 4684
rect 28215 4644 28488 4672
rect 29139 4644 29184 4672
rect 28215 4641 28227 4644
rect 28169 4635 28227 4641
rect 29178 4632 29184 4644
rect 29236 4632 29242 4684
rect 30650 4672 30656 4684
rect 30611 4644 30656 4672
rect 30650 4632 30656 4644
rect 30708 4632 30714 4684
rect 28077 4607 28135 4613
rect 28077 4573 28089 4607
rect 28123 4604 28135 4607
rect 28258 4604 28264 4616
rect 28123 4576 28264 4604
rect 28123 4573 28135 4576
rect 28077 4567 28135 4573
rect 28258 4564 28264 4576
rect 28316 4604 28322 4616
rect 28537 4607 28595 4613
rect 28537 4604 28549 4607
rect 28316 4576 28549 4604
rect 28316 4564 28322 4576
rect 28537 4573 28549 4576
rect 28583 4573 28595 4607
rect 28537 4567 28595 4573
rect 28997 4539 29055 4545
rect 28997 4536 29009 4539
rect 27908 4508 29009 4536
rect 28997 4505 29009 4508
rect 29043 4505 29055 4539
rect 28997 4499 29055 4505
rect 20496 4440 21864 4468
rect 25639 4471 25697 4477
rect 20496 4428 20502 4440
rect 25639 4437 25651 4471
rect 25685 4468 25697 4471
rect 26602 4468 26608 4480
rect 25685 4440 26608 4468
rect 25685 4437 25697 4440
rect 25639 4431 25697 4437
rect 26602 4428 26608 4440
rect 26660 4428 26666 4480
rect 26694 4428 26700 4480
rect 26752 4468 26758 4480
rect 28350 4468 28356 4480
rect 26752 4440 28356 4468
rect 26752 4428 26758 4440
rect 28350 4428 28356 4440
rect 28408 4428 28414 4480
rect 30466 4468 30472 4480
rect 30427 4440 30472 4468
rect 30466 4428 30472 4440
rect 30524 4428 30530 4480
rect 1104 4378 38824 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 38824 4378
rect 1104 4304 38824 4326
rect 16114 4224 16120 4276
rect 16172 4264 16178 4276
rect 16209 4267 16267 4273
rect 16209 4264 16221 4267
rect 16172 4236 16221 4264
rect 16172 4224 16178 4236
rect 16209 4233 16221 4236
rect 16255 4233 16267 4267
rect 16209 4227 16267 4233
rect 16574 4224 16580 4276
rect 16632 4264 16638 4276
rect 17770 4264 17776 4276
rect 16632 4236 17776 4264
rect 16632 4224 16638 4236
rect 17770 4224 17776 4236
rect 17828 4264 17834 4276
rect 19978 4264 19984 4276
rect 17828 4236 19984 4264
rect 17828 4224 17834 4236
rect 19978 4224 19984 4236
rect 20036 4224 20042 4276
rect 20152 4267 20210 4273
rect 20152 4233 20164 4267
rect 20198 4264 20210 4267
rect 22922 4264 22928 4276
rect 20198 4236 22928 4264
rect 20198 4233 20210 4236
rect 20152 4227 20210 4233
rect 22922 4224 22928 4236
rect 22980 4224 22986 4276
rect 25212 4267 25270 4273
rect 25212 4233 25224 4267
rect 25258 4264 25270 4267
rect 27430 4264 27436 4276
rect 25258 4236 27436 4264
rect 25258 4233 25270 4236
rect 25212 4227 25270 4233
rect 27430 4224 27436 4236
rect 27488 4224 27494 4276
rect 27798 4264 27804 4276
rect 27759 4236 27804 4264
rect 27798 4224 27804 4236
rect 27856 4224 27862 4276
rect 23106 4196 23112 4208
rect 17236 4168 17816 4196
rect 17236 4128 17264 4168
rect 14936 4100 17264 4128
rect 14936 4069 14964 4100
rect 17310 4088 17316 4140
rect 17368 4128 17374 4140
rect 17681 4131 17739 4137
rect 17681 4128 17693 4131
rect 17368 4100 17693 4128
rect 17368 4088 17374 4100
rect 17681 4097 17693 4100
rect 17727 4097 17739 4131
rect 17788 4128 17816 4168
rect 22204 4168 23112 4196
rect 18506 4128 18512 4140
rect 17788 4100 18512 4128
rect 17681 4091 17739 4097
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 18598 4088 18604 4140
rect 18656 4128 18662 4140
rect 22204 4128 22232 4168
rect 23106 4156 23112 4168
rect 23164 4156 23170 4208
rect 30466 4196 30472 4208
rect 26252 4168 30472 4196
rect 18656 4100 22232 4128
rect 18656 4088 18662 4100
rect 22278 4088 22284 4140
rect 22336 4128 22342 4140
rect 22649 4131 22707 4137
rect 22649 4128 22661 4131
rect 22336 4100 22661 4128
rect 22336 4088 22342 4100
rect 22649 4097 22661 4100
rect 22695 4097 22707 4131
rect 22649 4091 22707 4097
rect 24854 4088 24860 4140
rect 24912 4128 24918 4140
rect 26252 4128 26280 4168
rect 30466 4156 30472 4168
rect 30524 4156 30530 4208
rect 27614 4128 27620 4140
rect 24912 4100 26280 4128
rect 26344 4100 27620 4128
rect 24912 4088 24918 4100
rect 14921 4063 14979 4069
rect 14921 4029 14933 4063
rect 14967 4029 14979 4063
rect 14921 4023 14979 4029
rect 15565 4063 15623 4069
rect 15565 4029 15577 4063
rect 15611 4060 15623 4063
rect 16114 4060 16120 4072
rect 15611 4032 16120 4060
rect 15611 4029 15623 4032
rect 15565 4023 15623 4029
rect 16114 4020 16120 4032
rect 16172 4020 16178 4072
rect 16390 4060 16396 4072
rect 16351 4032 16396 4060
rect 16390 4020 16396 4032
rect 16448 4020 16454 4072
rect 19426 4020 19432 4072
rect 19484 4060 19490 4072
rect 19889 4063 19947 4069
rect 19889 4060 19901 4063
rect 19484 4032 19901 4060
rect 19484 4020 19490 4032
rect 19889 4029 19901 4032
rect 19935 4029 19947 4063
rect 19889 4023 19947 4029
rect 24397 4063 24455 4069
rect 24397 4029 24409 4063
rect 24443 4060 24455 4063
rect 24949 4063 25007 4069
rect 24949 4060 24961 4063
rect 24443 4032 24961 4060
rect 24443 4029 24455 4032
rect 24397 4023 24455 4029
rect 24949 4029 24961 4032
rect 24995 4029 25007 4063
rect 26344 4046 26372 4100
rect 27614 4088 27620 4100
rect 27672 4088 27678 4140
rect 27890 4088 27896 4140
rect 27948 4128 27954 4140
rect 28353 4131 28411 4137
rect 28353 4128 28365 4131
rect 27948 4100 28365 4128
rect 27948 4088 27954 4100
rect 28092 4069 28120 4100
rect 28353 4097 28365 4100
rect 28399 4097 28411 4131
rect 30650 4128 30656 4140
rect 28353 4091 28411 4097
rect 29748 4100 30656 4128
rect 27985 4063 28043 4069
rect 24949 4023 25007 4029
rect 27985 4029 27997 4063
rect 28031 4029 28043 4063
rect 27985 4023 28043 4029
rect 28077 4063 28135 4069
rect 28077 4029 28089 4063
rect 28123 4029 28135 4063
rect 28077 4023 28135 4029
rect 17954 3992 17960 4004
rect 15120 3964 17816 3992
rect 17915 3964 17960 3992
rect 15120 3933 15148 3964
rect 15105 3927 15163 3933
rect 15105 3893 15117 3927
rect 15151 3893 15163 3927
rect 15105 3887 15163 3893
rect 15749 3927 15807 3933
rect 15749 3893 15761 3927
rect 15795 3924 15807 3927
rect 17678 3924 17684 3936
rect 15795 3896 17684 3924
rect 15795 3893 15807 3896
rect 15749 3887 15807 3893
rect 17678 3884 17684 3896
rect 17736 3884 17742 3936
rect 17788 3924 17816 3964
rect 17954 3952 17960 3964
rect 18012 3952 18018 4004
rect 19242 3992 19248 4004
rect 19182 3964 19248 3992
rect 19242 3952 19248 3964
rect 19300 3952 19306 4004
rect 20438 3992 20444 4004
rect 19352 3964 20444 3992
rect 19352 3924 19380 3964
rect 20438 3952 20444 3964
rect 20496 3952 20502 4004
rect 22830 3992 22836 4004
rect 21390 3964 22836 3992
rect 22830 3952 22836 3964
rect 22888 3952 22894 4004
rect 23658 3952 23664 4004
rect 23716 3952 23722 4004
rect 24121 3995 24179 4001
rect 24121 3961 24133 3995
rect 24167 3992 24179 3995
rect 24210 3992 24216 4004
rect 24167 3964 24216 3992
rect 24167 3961 24179 3964
rect 24121 3955 24179 3961
rect 24210 3952 24216 3964
rect 24268 3952 24274 4004
rect 24964 3992 24992 4023
rect 25222 3992 25228 4004
rect 24964 3964 25228 3992
rect 25222 3952 25228 3964
rect 25280 3952 25286 4004
rect 27890 3992 27896 4004
rect 26528 3964 27896 3992
rect 17788 3896 19380 3924
rect 19429 3927 19487 3933
rect 19429 3893 19441 3927
rect 19475 3924 19487 3927
rect 21450 3924 21456 3936
rect 19475 3896 21456 3924
rect 19475 3893 19487 3896
rect 19429 3887 19487 3893
rect 21450 3884 21456 3896
rect 21508 3884 21514 3936
rect 21637 3927 21695 3933
rect 21637 3893 21649 3927
rect 21683 3924 21695 3927
rect 22462 3924 22468 3936
rect 21683 3896 22468 3924
rect 21683 3893 21695 3896
rect 21637 3887 21695 3893
rect 22462 3884 22468 3896
rect 22520 3884 22526 3936
rect 22646 3884 22652 3936
rect 22704 3924 22710 3936
rect 26528 3924 26556 3964
rect 27890 3952 27896 3964
rect 27948 3952 27954 4004
rect 28000 3992 28028 4023
rect 28166 4020 28172 4072
rect 28224 4060 28230 4072
rect 29089 4063 29147 4069
rect 29089 4060 29101 4063
rect 28224 4032 29101 4060
rect 28224 4020 28230 4032
rect 29089 4029 29101 4032
rect 29135 4060 29147 4063
rect 29362 4060 29368 4072
rect 29135 4032 29368 4060
rect 29135 4029 29147 4032
rect 29089 4023 29147 4029
rect 29362 4020 29368 4032
rect 29420 4020 29426 4072
rect 29748 4069 29776 4100
rect 30650 4088 30656 4100
rect 30708 4088 30714 4140
rect 29733 4063 29791 4069
rect 29733 4029 29745 4063
rect 29779 4029 29791 4063
rect 29733 4023 29791 4029
rect 30193 4063 30251 4069
rect 30193 4029 30205 4063
rect 30239 4029 30251 4063
rect 30193 4023 30251 4029
rect 28258 3992 28264 4004
rect 28000 3964 28264 3992
rect 28258 3952 28264 3964
rect 28316 3992 28322 4004
rect 28445 3995 28503 4001
rect 28445 3992 28457 3995
rect 28316 3964 28457 3992
rect 28316 3952 28322 3964
rect 28445 3961 28457 3964
rect 28491 3961 28503 3995
rect 30208 3992 30236 4023
rect 28445 3955 28503 3961
rect 28552 3964 30236 3992
rect 26694 3924 26700 3936
rect 22704 3896 26556 3924
rect 26607 3896 26700 3924
rect 22704 3884 22710 3896
rect 26694 3884 26700 3896
rect 26752 3924 26758 3936
rect 28552 3924 28580 3964
rect 26752 3896 28580 3924
rect 26752 3884 26758 3896
rect 28626 3884 28632 3936
rect 28684 3924 28690 3936
rect 28905 3927 28963 3933
rect 28905 3924 28917 3927
rect 28684 3896 28917 3924
rect 28684 3884 28690 3896
rect 28905 3893 28917 3896
rect 28951 3893 28963 3927
rect 28905 3887 28963 3893
rect 28994 3884 29000 3936
rect 29052 3924 29058 3936
rect 29549 3927 29607 3933
rect 29549 3924 29561 3927
rect 29052 3896 29561 3924
rect 29052 3884 29058 3896
rect 29549 3893 29561 3896
rect 29595 3893 29607 3927
rect 29549 3887 29607 3893
rect 29638 3884 29644 3936
rect 29696 3924 29702 3936
rect 30285 3927 30343 3933
rect 30285 3924 30297 3927
rect 29696 3896 30297 3924
rect 29696 3884 29702 3896
rect 30285 3893 30297 3896
rect 30331 3893 30343 3927
rect 30285 3887 30343 3893
rect 1104 3834 38824 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 38824 3834
rect 1104 3760 38824 3782
rect 16853 3723 16911 3729
rect 16853 3689 16865 3723
rect 16899 3720 16911 3723
rect 19061 3723 19119 3729
rect 16899 3692 19012 3720
rect 16899 3689 16911 3692
rect 16853 3683 16911 3689
rect 16574 3652 16580 3664
rect 16040 3624 16580 3652
rect 15746 3544 15752 3596
rect 15804 3584 15810 3596
rect 16040 3593 16068 3624
rect 16574 3612 16580 3624
rect 16632 3612 16638 3664
rect 17586 3652 17592 3664
rect 17547 3624 17592 3652
rect 17586 3612 17592 3624
rect 17644 3612 17650 3664
rect 18598 3612 18604 3664
rect 18656 3612 18662 3664
rect 18984 3652 19012 3692
rect 19061 3689 19073 3723
rect 19107 3720 19119 3723
rect 19107 3692 24164 3720
rect 19107 3689 19119 3692
rect 19061 3683 19119 3689
rect 18984 3624 20654 3652
rect 22370 3612 22376 3664
rect 22428 3652 22434 3664
rect 22833 3655 22891 3661
rect 22833 3652 22845 3655
rect 22428 3624 22845 3652
rect 22428 3612 22434 3624
rect 22833 3621 22845 3624
rect 22879 3621 22891 3655
rect 24136 3652 24164 3692
rect 24210 3680 24216 3732
rect 24268 3720 24274 3732
rect 24305 3723 24363 3729
rect 24305 3720 24317 3723
rect 24268 3692 24317 3720
rect 24268 3680 24274 3692
rect 24305 3689 24317 3692
rect 24351 3689 24363 3723
rect 24305 3683 24363 3689
rect 24578 3680 24584 3732
rect 24636 3720 24642 3732
rect 26973 3723 27031 3729
rect 24636 3692 26832 3720
rect 24636 3680 24642 3692
rect 25501 3655 25559 3661
rect 25501 3652 25513 3655
rect 24136 3624 25513 3652
rect 22833 3615 22891 3621
rect 25501 3621 25513 3624
rect 25547 3621 25559 3655
rect 26804 3652 26832 3692
rect 26973 3689 26985 3723
rect 27019 3720 27031 3723
rect 27062 3720 27068 3732
rect 27019 3692 27068 3720
rect 27019 3689 27031 3692
rect 26973 3683 27031 3689
rect 27062 3680 27068 3692
rect 27120 3680 27126 3732
rect 27614 3680 27620 3732
rect 27672 3720 27678 3732
rect 29365 3723 29423 3729
rect 29365 3720 29377 3723
rect 27672 3692 29377 3720
rect 27672 3680 27678 3692
rect 29365 3689 29377 3692
rect 29411 3689 29423 3723
rect 29365 3683 29423 3689
rect 28994 3652 29000 3664
rect 26804 3624 29000 3652
rect 25501 3615 25559 3621
rect 28994 3612 29000 3624
rect 29052 3612 29058 3664
rect 16025 3587 16083 3593
rect 16025 3584 16037 3587
rect 15804 3556 16037 3584
rect 15804 3544 15810 3556
rect 16025 3553 16037 3556
rect 16071 3553 16083 3587
rect 16025 3547 16083 3553
rect 16114 3544 16120 3596
rect 16172 3584 16178 3596
rect 16669 3587 16727 3593
rect 16669 3584 16681 3587
rect 16172 3556 16681 3584
rect 16172 3544 16178 3556
rect 16669 3553 16681 3556
rect 16715 3553 16727 3587
rect 17310 3584 17316 3596
rect 17271 3556 17316 3584
rect 16669 3547 16727 3553
rect 16684 3448 16712 3547
rect 17310 3544 17316 3556
rect 17368 3544 17374 3596
rect 22097 3587 22155 3593
rect 22097 3553 22109 3587
rect 22143 3584 22155 3587
rect 22186 3584 22192 3596
rect 22143 3556 22192 3584
rect 22143 3553 22155 3556
rect 22097 3547 22155 3553
rect 22186 3544 22192 3556
rect 22244 3584 22250 3596
rect 22554 3584 22560 3596
rect 22244 3556 22560 3584
rect 22244 3544 22250 3556
rect 22554 3544 22560 3556
rect 22612 3544 22618 3596
rect 24854 3584 24860 3596
rect 23966 3556 24860 3584
rect 24854 3544 24860 3556
rect 24912 3544 24918 3596
rect 25222 3584 25228 3596
rect 25183 3556 25228 3584
rect 25222 3544 25228 3556
rect 25280 3544 25286 3596
rect 27246 3584 27252 3596
rect 26634 3556 27252 3584
rect 27246 3544 27252 3556
rect 27304 3544 27310 3596
rect 27338 3544 27344 3596
rect 27396 3584 27402 3596
rect 27433 3587 27491 3593
rect 27433 3584 27445 3587
rect 27396 3556 27445 3584
rect 27396 3544 27402 3556
rect 27433 3553 27445 3556
rect 27479 3553 27491 3587
rect 27433 3547 27491 3553
rect 28166 3544 28172 3596
rect 28224 3584 28230 3596
rect 28261 3587 28319 3593
rect 28261 3584 28273 3587
rect 28224 3556 28273 3584
rect 28224 3544 28230 3556
rect 28261 3553 28273 3556
rect 28307 3553 28319 3587
rect 28261 3547 28319 3553
rect 28534 3544 28540 3596
rect 28592 3584 28598 3596
rect 28902 3584 28908 3596
rect 28592 3556 28908 3584
rect 28592 3544 28598 3556
rect 28902 3544 28908 3556
rect 28960 3544 28966 3596
rect 29546 3584 29552 3596
rect 29507 3556 29552 3584
rect 29546 3544 29552 3556
rect 29604 3584 29610 3596
rect 31386 3584 31392 3596
rect 29604 3556 31392 3584
rect 29604 3544 29610 3556
rect 31386 3544 31392 3556
rect 31444 3544 31450 3596
rect 17420 3488 18644 3516
rect 17420 3448 17448 3488
rect 16684 3420 17448 3448
rect 18616 3448 18644 3488
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 21821 3519 21879 3525
rect 21821 3516 21833 3519
rect 19484 3488 21833 3516
rect 19484 3476 19490 3488
rect 21821 3485 21833 3488
rect 21867 3485 21879 3519
rect 26786 3516 26792 3528
rect 21821 3479 21879 3485
rect 22066 3488 23888 3516
rect 18616 3420 20484 3448
rect 16117 3383 16175 3389
rect 16117 3349 16129 3383
rect 16163 3380 16175 3383
rect 18046 3380 18052 3392
rect 16163 3352 18052 3380
rect 16163 3349 16175 3352
rect 16117 3343 16175 3349
rect 18046 3340 18052 3352
rect 18104 3340 18110 3392
rect 20346 3380 20352 3392
rect 20307 3352 20352 3380
rect 20346 3340 20352 3352
rect 20404 3340 20410 3392
rect 20456 3380 20484 3420
rect 22066 3380 22094 3488
rect 23860 3448 23888 3488
rect 25332 3488 26792 3516
rect 25332 3448 25360 3488
rect 26786 3476 26792 3488
rect 26844 3476 26850 3528
rect 27890 3476 27896 3528
rect 27948 3516 27954 3528
rect 27948 3488 28120 3516
rect 27948 3476 27954 3488
rect 23860 3420 25360 3448
rect 27617 3451 27675 3457
rect 27617 3417 27629 3451
rect 27663 3448 27675 3451
rect 27982 3448 27988 3460
rect 27663 3420 27988 3448
rect 27663 3417 27675 3420
rect 27617 3411 27675 3417
rect 27982 3408 27988 3420
rect 28040 3408 28046 3460
rect 28092 3457 28120 3488
rect 28350 3476 28356 3528
rect 28408 3516 28414 3528
rect 28408 3488 31754 3516
rect 28408 3476 28414 3488
rect 31726 3460 31754 3488
rect 28077 3451 28135 3457
rect 28077 3417 28089 3451
rect 28123 3417 28135 3451
rect 31726 3420 31760 3460
rect 28077 3411 28135 3417
rect 31754 3408 31760 3420
rect 31812 3408 31818 3460
rect 20456 3352 22094 3380
rect 22830 3340 22836 3392
rect 22888 3380 22894 3392
rect 28721 3383 28779 3389
rect 28721 3380 28733 3383
rect 22888 3352 28733 3380
rect 22888 3340 22894 3352
rect 28721 3349 28733 3352
rect 28767 3349 28779 3383
rect 28721 3343 28779 3349
rect 1104 3290 38824 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 38824 3290
rect 1104 3216 38824 3238
rect 17770 3136 17776 3188
rect 17828 3176 17834 3188
rect 17865 3179 17923 3185
rect 17865 3176 17877 3179
rect 17828 3148 17877 3176
rect 17828 3136 17834 3148
rect 17865 3145 17877 3148
rect 17911 3145 17923 3179
rect 17865 3139 17923 3145
rect 17954 3136 17960 3188
rect 18012 3176 18018 3188
rect 18325 3179 18383 3185
rect 18325 3176 18337 3179
rect 18012 3148 18337 3176
rect 18012 3136 18018 3148
rect 18325 3145 18337 3148
rect 18371 3145 18383 3179
rect 19426 3176 19432 3188
rect 19387 3148 19432 3176
rect 18325 3139 18383 3145
rect 19426 3136 19432 3148
rect 19484 3136 19490 3188
rect 19889 3179 19947 3185
rect 19889 3145 19901 3179
rect 19935 3176 19947 3179
rect 20070 3176 20076 3188
rect 19935 3148 20076 3176
rect 19935 3145 19947 3148
rect 19889 3139 19947 3145
rect 20070 3136 20076 3148
rect 20128 3136 20134 3188
rect 21174 3136 21180 3188
rect 21232 3176 21238 3188
rect 24305 3179 24363 3185
rect 24305 3176 24317 3179
rect 21232 3148 24317 3176
rect 21232 3136 21238 3148
rect 24305 3145 24317 3148
rect 24351 3145 24363 3179
rect 24305 3139 24363 3145
rect 26145 3179 26203 3185
rect 26145 3145 26157 3179
rect 26191 3176 26203 3179
rect 26326 3176 26332 3188
rect 26191 3148 26332 3176
rect 26191 3145 26203 3148
rect 26145 3139 26203 3145
rect 26326 3136 26332 3148
rect 26384 3136 26390 3188
rect 26602 3176 26608 3188
rect 26563 3148 26608 3176
rect 26602 3136 26608 3148
rect 26660 3176 26666 3188
rect 26878 3176 26884 3188
rect 26660 3148 26884 3176
rect 26660 3136 26666 3148
rect 26878 3136 26884 3148
rect 26936 3136 26942 3188
rect 26970 3136 26976 3188
rect 27028 3176 27034 3188
rect 29178 3176 29184 3188
rect 27028 3148 29184 3176
rect 27028 3136 27034 3148
rect 29178 3136 29184 3148
rect 29236 3136 29242 3188
rect 17494 3068 17500 3120
rect 17552 3108 17558 3120
rect 25593 3111 25651 3117
rect 17552 3080 19380 3108
rect 17552 3068 17558 3080
rect 19245 3043 19303 3049
rect 19245 3040 19257 3043
rect 18064 3012 18276 3040
rect 18064 2984 18092 3012
rect 15102 2932 15108 2984
rect 15160 2972 15166 2984
rect 17773 2975 17831 2981
rect 17773 2972 17785 2975
rect 15160 2944 17785 2972
rect 15160 2932 15166 2944
rect 17773 2941 17785 2944
rect 17819 2941 17831 2975
rect 18046 2972 18052 2984
rect 18007 2944 18052 2972
rect 17773 2935 17831 2941
rect 18046 2932 18052 2944
rect 18104 2932 18110 2984
rect 18141 2975 18199 2981
rect 18141 2941 18153 2975
rect 18187 2941 18199 2975
rect 18248 2972 18276 3012
rect 18800 3012 19257 3040
rect 18690 2972 18696 2984
rect 18248 2944 18696 2972
rect 18141 2935 18199 2941
rect 16482 2864 16488 2916
rect 16540 2904 16546 2916
rect 18156 2904 18184 2935
rect 18690 2932 18696 2944
rect 18748 2972 18754 2984
rect 18800 2981 18828 3012
rect 19245 3009 19257 3012
rect 19291 3009 19303 3043
rect 19245 3003 19303 3009
rect 18785 2975 18843 2981
rect 18785 2972 18797 2975
rect 18748 2944 18797 2972
rect 18748 2932 18754 2944
rect 18785 2941 18797 2944
rect 18831 2941 18843 2975
rect 18785 2935 18843 2941
rect 18877 2975 18935 2981
rect 18877 2941 18889 2975
rect 18923 2972 18935 2975
rect 19150 2972 19156 2984
rect 18923 2944 19156 2972
rect 18923 2941 18935 2944
rect 18877 2935 18935 2941
rect 19150 2932 19156 2944
rect 19208 2932 19214 2984
rect 19352 2972 19380 3080
rect 25593 3077 25605 3111
rect 25639 3108 25651 3111
rect 26234 3108 26240 3120
rect 25639 3080 26240 3108
rect 25639 3077 25651 3080
rect 25593 3071 25651 3077
rect 26234 3068 26240 3080
rect 26292 3068 26298 3120
rect 27062 3068 27068 3120
rect 27120 3108 27126 3120
rect 29089 3111 29147 3117
rect 29089 3108 29101 3111
rect 27120 3080 29101 3108
rect 27120 3068 27126 3080
rect 29089 3077 29101 3080
rect 29135 3077 29147 3111
rect 30193 3111 30251 3117
rect 30193 3108 30205 3111
rect 29089 3071 29147 3077
rect 29748 3080 30205 3108
rect 20622 3000 20628 3052
rect 20680 3040 20686 3052
rect 21361 3043 21419 3049
rect 21361 3040 21373 3043
rect 20680 3012 21373 3040
rect 20680 3000 20686 3012
rect 21361 3009 21373 3012
rect 21407 3009 21419 3043
rect 21361 3003 21419 3009
rect 21637 3043 21695 3049
rect 21637 3009 21649 3043
rect 21683 3040 21695 3043
rect 22186 3040 22192 3052
rect 21683 3012 22192 3040
rect 21683 3009 21695 3012
rect 21637 3003 21695 3009
rect 22186 3000 22192 3012
rect 22244 3000 22250 3052
rect 22462 3000 22468 3052
rect 22520 3040 22526 3052
rect 22833 3043 22891 3049
rect 22833 3040 22845 3043
rect 22520 3012 22845 3040
rect 22520 3000 22526 3012
rect 22833 3009 22845 3012
rect 22879 3009 22891 3043
rect 29638 3040 29644 3052
rect 22833 3003 22891 3009
rect 26344 3012 29644 3040
rect 22204 2972 22232 3000
rect 22557 2975 22615 2981
rect 22557 2972 22569 2975
rect 19352 2944 20286 2972
rect 22204 2944 22569 2972
rect 22557 2941 22569 2944
rect 22603 2941 22615 2975
rect 22557 2935 22615 2941
rect 24670 2932 24676 2984
rect 24728 2972 24734 2984
rect 24765 2975 24823 2981
rect 24765 2972 24777 2975
rect 24728 2944 24777 2972
rect 24728 2932 24734 2944
rect 24765 2941 24777 2944
rect 24811 2941 24823 2975
rect 25409 2975 25467 2981
rect 25409 2972 25421 2975
rect 24765 2935 24823 2941
rect 24964 2944 25421 2972
rect 24578 2904 24584 2916
rect 16540 2876 18184 2904
rect 24058 2876 24584 2904
rect 16540 2864 16546 2876
rect 24578 2864 24584 2876
rect 24636 2864 24642 2916
rect 11146 2836 11152 2848
rect 11107 2808 11152 2836
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 16390 2796 16396 2848
rect 16448 2836 16454 2848
rect 24964 2845 24992 2944
rect 25409 2941 25421 2944
rect 25455 2972 25467 2975
rect 25774 2972 25780 2984
rect 25455 2944 25780 2972
rect 25455 2941 25467 2944
rect 25409 2935 25467 2941
rect 25774 2932 25780 2944
rect 25832 2932 25838 2984
rect 26344 2981 26372 3012
rect 29638 3000 29644 3012
rect 29696 3000 29702 3052
rect 29748 3049 29776 3080
rect 30193 3077 30205 3080
rect 30239 3077 30251 3111
rect 30193 3071 30251 3077
rect 29733 3043 29791 3049
rect 29733 3009 29745 3043
rect 29779 3009 29791 3043
rect 29733 3003 29791 3009
rect 26329 2975 26387 2981
rect 26329 2941 26341 2975
rect 26375 2941 26387 2975
rect 26329 2935 26387 2941
rect 26421 2975 26479 2981
rect 26421 2941 26433 2975
rect 26467 2941 26479 2975
rect 26694 2972 26700 2984
rect 26655 2944 26700 2972
rect 26421 2935 26479 2941
rect 26436 2904 26464 2935
rect 26694 2932 26700 2944
rect 26752 2932 26758 2984
rect 27985 2975 28043 2981
rect 27985 2941 27997 2975
rect 28031 2972 28043 2975
rect 28350 2972 28356 2984
rect 28031 2944 28356 2972
rect 28031 2941 28043 2944
rect 27985 2935 28043 2941
rect 28350 2932 28356 2944
rect 28408 2932 28414 2984
rect 28629 2975 28687 2981
rect 28629 2941 28641 2975
rect 28675 2972 28687 2975
rect 29546 2972 29552 2984
rect 28675 2944 29552 2972
rect 28675 2941 28687 2944
rect 28629 2935 28687 2941
rect 29546 2932 29552 2944
rect 29604 2932 29610 2984
rect 30377 2975 30435 2981
rect 30377 2941 30389 2975
rect 30423 2941 30435 2975
rect 30377 2935 30435 2941
rect 28258 2904 28264 2916
rect 26436 2876 28264 2904
rect 28258 2864 28264 2876
rect 28316 2864 28322 2916
rect 28718 2864 28724 2916
rect 28776 2904 28782 2916
rect 30392 2904 30420 2935
rect 28776 2876 30420 2904
rect 28776 2864 28782 2876
rect 24949 2839 25007 2845
rect 24949 2836 24961 2839
rect 16448 2808 24961 2836
rect 16448 2796 16454 2808
rect 24949 2805 24961 2808
rect 24995 2805 25007 2839
rect 24949 2799 25007 2805
rect 25038 2796 25044 2848
rect 25096 2836 25102 2848
rect 27801 2839 27859 2845
rect 27801 2836 27813 2839
rect 25096 2808 27813 2836
rect 25096 2796 25102 2808
rect 27801 2805 27813 2808
rect 27847 2805 27859 2839
rect 28442 2836 28448 2848
rect 28403 2808 28448 2836
rect 27801 2799 27859 2805
rect 28442 2796 28448 2808
rect 28500 2796 28506 2848
rect 1104 2746 38824 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 38824 2746
rect 1104 2672 38824 2694
rect 19337 2635 19395 2641
rect 19337 2601 19349 2635
rect 19383 2632 19395 2635
rect 20714 2632 20720 2644
rect 19383 2604 20720 2632
rect 19383 2601 19395 2604
rect 19337 2595 19395 2601
rect 20714 2592 20720 2604
rect 20772 2592 20778 2644
rect 22922 2632 22928 2644
rect 22883 2604 22928 2632
rect 22922 2592 22928 2604
rect 22980 2592 22986 2644
rect 23106 2592 23112 2644
rect 23164 2632 23170 2644
rect 25593 2635 25651 2641
rect 25593 2632 25605 2635
rect 23164 2604 25605 2632
rect 23164 2592 23170 2604
rect 25593 2601 25605 2604
rect 25639 2601 25651 2635
rect 25593 2595 25651 2601
rect 25774 2592 25780 2644
rect 25832 2632 25838 2644
rect 26237 2635 26295 2641
rect 25832 2604 25912 2632
rect 25832 2592 25838 2604
rect 11146 2524 11152 2576
rect 11204 2564 11210 2576
rect 11241 2567 11299 2573
rect 11241 2564 11253 2567
rect 11204 2536 11253 2564
rect 11204 2524 11210 2536
rect 11241 2533 11253 2536
rect 11287 2533 11299 2567
rect 15746 2564 15752 2576
rect 15707 2536 15752 2564
rect 11241 2527 11299 2533
rect 15746 2524 15752 2536
rect 15804 2524 15810 2576
rect 18690 2564 18696 2576
rect 18651 2536 18696 2564
rect 18690 2524 18696 2536
rect 18748 2524 18754 2576
rect 21082 2524 21088 2576
rect 21140 2524 21146 2576
rect 21450 2524 21456 2576
rect 21508 2564 21514 2576
rect 21729 2567 21787 2573
rect 21729 2564 21741 2567
rect 21508 2536 21741 2564
rect 21508 2524 21514 2536
rect 21729 2533 21741 2536
rect 21775 2533 21787 2567
rect 25038 2564 25044 2576
rect 23966 2536 25044 2564
rect 21729 2527 21787 2533
rect 25038 2524 25044 2536
rect 25096 2524 25102 2576
rect 25884 2564 25912 2604
rect 26237 2601 26249 2635
rect 26283 2632 26295 2635
rect 26602 2632 26608 2644
rect 26283 2604 26608 2632
rect 26283 2601 26295 2604
rect 26237 2595 26295 2601
rect 26602 2592 26608 2604
rect 26660 2592 26666 2644
rect 26878 2592 26884 2644
rect 26936 2632 26942 2644
rect 26936 2604 27108 2632
rect 26936 2592 26942 2604
rect 26970 2564 26976 2576
rect 25884 2536 26976 2564
rect 2409 2499 2467 2505
rect 2409 2465 2421 2499
rect 2455 2496 2467 2499
rect 2961 2499 3019 2505
rect 2961 2496 2973 2499
rect 2455 2468 2973 2496
rect 2455 2465 2467 2468
rect 2409 2459 2467 2465
rect 2961 2465 2973 2468
rect 3007 2465 3019 2499
rect 2961 2459 3019 2465
rect 16669 2499 16727 2505
rect 16669 2465 16681 2499
rect 16715 2496 16727 2499
rect 18049 2499 18107 2505
rect 18049 2496 18061 2499
rect 16715 2468 18061 2496
rect 16715 2465 16727 2468
rect 16669 2459 16727 2465
rect 18049 2465 18061 2468
rect 18095 2465 18107 2499
rect 18049 2459 18107 2465
rect 18708 2428 18736 2524
rect 18785 2499 18843 2505
rect 18785 2465 18797 2499
rect 18831 2496 18843 2499
rect 19061 2499 19119 2505
rect 19061 2496 19073 2499
rect 18831 2468 19073 2496
rect 18831 2465 18843 2468
rect 18785 2459 18843 2465
rect 19061 2465 19073 2468
rect 19107 2496 19119 2499
rect 20346 2496 20352 2508
rect 19107 2468 20352 2496
rect 19107 2465 19119 2468
rect 19061 2459 19119 2465
rect 20346 2456 20352 2468
rect 20404 2456 20410 2508
rect 22005 2499 22063 2505
rect 22005 2465 22017 2499
rect 22051 2496 22063 2499
rect 22278 2496 22284 2508
rect 22051 2468 22284 2496
rect 22051 2465 22063 2468
rect 22005 2459 22063 2465
rect 22278 2456 22284 2468
rect 22336 2456 22342 2508
rect 24673 2499 24731 2505
rect 24673 2465 24685 2499
rect 24719 2496 24731 2499
rect 25222 2496 25228 2508
rect 24719 2468 25228 2496
rect 24719 2465 24731 2468
rect 24673 2459 24731 2465
rect 25222 2456 25228 2468
rect 25280 2456 25286 2508
rect 25777 2499 25835 2505
rect 25777 2465 25789 2499
rect 25823 2496 25835 2499
rect 25884 2496 25912 2536
rect 26970 2524 26976 2536
rect 27028 2524 27034 2576
rect 27080 2564 27108 2604
rect 28258 2592 28264 2644
rect 28316 2632 28322 2644
rect 28353 2635 28411 2641
rect 28353 2632 28365 2635
rect 28316 2604 28365 2632
rect 28316 2592 28322 2604
rect 28353 2601 28365 2604
rect 28399 2601 28411 2635
rect 28353 2595 28411 2601
rect 33781 2567 33839 2573
rect 33781 2564 33793 2567
rect 27080 2536 33793 2564
rect 25823 2468 25912 2496
rect 26421 2499 26479 2505
rect 25823 2465 25835 2468
rect 25777 2459 25835 2465
rect 26421 2465 26433 2499
rect 26467 2465 26479 2499
rect 26421 2459 26479 2465
rect 19153 2431 19211 2437
rect 19153 2428 19165 2431
rect 18708 2400 19165 2428
rect 19153 2397 19165 2400
rect 19199 2397 19211 2431
rect 20254 2428 20260 2440
rect 20215 2400 20260 2428
rect 19153 2391 19211 2397
rect 20254 2388 20260 2400
rect 20312 2388 20318 2440
rect 24397 2431 24455 2437
rect 24397 2397 24409 2431
rect 24443 2428 24455 2431
rect 26436 2428 26464 2459
rect 26786 2456 26792 2508
rect 26844 2496 26850 2508
rect 27065 2499 27123 2505
rect 27065 2496 27077 2499
rect 26844 2468 27077 2496
rect 26844 2456 26850 2468
rect 27065 2465 27077 2468
rect 27111 2496 27123 2499
rect 28350 2496 28356 2508
rect 27111 2468 28356 2496
rect 27111 2465 27123 2468
rect 27065 2459 27123 2465
rect 28350 2456 28356 2468
rect 28408 2456 28414 2508
rect 28460 2505 28488 2536
rect 33781 2533 33793 2536
rect 33827 2533 33839 2567
rect 33781 2527 33839 2533
rect 28445 2499 28503 2505
rect 28445 2465 28457 2499
rect 28491 2465 28503 2499
rect 28445 2459 28503 2465
rect 29089 2499 29147 2505
rect 29089 2465 29101 2499
rect 29135 2496 29147 2499
rect 29641 2499 29699 2505
rect 29641 2496 29653 2499
rect 29135 2468 29653 2496
rect 29135 2465 29147 2468
rect 29089 2459 29147 2465
rect 29641 2465 29653 2468
rect 29687 2465 29699 2499
rect 29641 2459 29699 2465
rect 37277 2499 37335 2505
rect 37277 2465 37289 2499
rect 37323 2496 37335 2499
rect 37921 2499 37979 2505
rect 37921 2496 37933 2499
rect 37323 2468 37933 2496
rect 37323 2465 37335 2468
rect 37277 2459 37335 2465
rect 37921 2465 37933 2468
rect 37967 2465 37979 2499
rect 37921 2459 37979 2465
rect 28166 2428 28172 2440
rect 24443 2400 26372 2428
rect 26436 2400 28172 2428
rect 24443 2397 24455 2400
rect 24397 2391 24455 2397
rect 2222 2360 2228 2372
rect 2183 2332 2228 2360
rect 2222 2320 2228 2332
rect 2280 2320 2286 2372
rect 11054 2360 11060 2372
rect 11015 2332 11060 2360
rect 11054 2320 11060 2332
rect 11112 2320 11118 2372
rect 15562 2360 15568 2372
rect 15523 2332 15568 2360
rect 15562 2320 15568 2332
rect 15620 2320 15626 2372
rect 18233 2363 18291 2369
rect 18233 2329 18245 2363
rect 18279 2360 18291 2363
rect 19978 2360 19984 2372
rect 18279 2332 19984 2360
rect 18279 2329 18291 2332
rect 18233 2323 18291 2329
rect 19978 2320 19984 2332
rect 20036 2320 20042 2372
rect 26344 2360 26372 2400
rect 28166 2388 28172 2400
rect 28224 2388 28230 2440
rect 27062 2360 27068 2372
rect 26344 2332 27068 2360
rect 27062 2320 27068 2332
rect 27120 2320 27126 2372
rect 28902 2360 28908 2372
rect 28863 2332 28908 2360
rect 28902 2320 28908 2332
rect 28960 2320 28966 2372
rect 33318 2320 33324 2372
rect 33376 2360 33382 2372
rect 33597 2363 33655 2369
rect 33597 2360 33609 2363
rect 33376 2332 33609 2360
rect 33376 2320 33382 2332
rect 33597 2329 33609 2332
rect 33643 2329 33655 2363
rect 37734 2360 37740 2372
rect 37695 2332 37740 2360
rect 33597 2323 33655 2329
rect 37734 2320 37740 2332
rect 37792 2320 37798 2372
rect 22094 2252 22100 2304
rect 22152 2292 22158 2304
rect 26881 2295 26939 2301
rect 26881 2292 26893 2295
rect 22152 2264 26893 2292
rect 22152 2252 22158 2264
rect 26881 2261 26893 2264
rect 26927 2261 26939 2295
rect 26881 2255 26939 2261
rect 1104 2202 38824 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 38824 2202
rect 1104 2128 38824 2150
rect 24394 960 24400 1012
rect 24452 1000 24458 1012
rect 28718 1000 28724 1012
rect 24452 972 28724 1000
rect 24452 960 24458 972
rect 28718 960 28724 972
rect 28776 960 28782 1012
<< via1 >>
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 20812 37272 20864 37324
rect 20444 37247 20496 37256
rect 20444 37213 20453 37247
rect 20453 37213 20487 37247
rect 20487 37213 20496 37247
rect 20444 37204 20496 37213
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 20444 36907 20496 36916
rect 20444 36873 20453 36907
rect 20453 36873 20487 36907
rect 20487 36873 20496 36907
rect 20444 36864 20496 36873
rect 19984 36660 20036 36712
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 19984 21496 20036 21548
rect 19064 21471 19116 21480
rect 19064 21437 19073 21471
rect 19073 21437 19107 21471
rect 19107 21437 19116 21471
rect 19064 21428 19116 21437
rect 20812 21360 20864 21412
rect 20352 21292 20404 21344
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 20812 21088 20864 21140
rect 19064 20995 19116 21004
rect 19064 20961 19073 20995
rect 19073 20961 19107 20995
rect 19107 20961 19116 20995
rect 19064 20952 19116 20961
rect 19984 20995 20036 21004
rect 19984 20961 19993 20995
rect 19993 20961 20027 20995
rect 20027 20961 20036 20995
rect 19984 20952 20036 20961
rect 20352 20995 20404 21004
rect 20352 20961 20361 20995
rect 20361 20961 20395 20995
rect 20395 20961 20404 20995
rect 20352 20952 20404 20961
rect 20904 20748 20956 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 19984 20408 20036 20460
rect 20904 20408 20956 20460
rect 20812 20272 20864 20324
rect 21640 20204 21692 20256
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 20812 19932 20864 19984
rect 21640 19907 21692 19916
rect 21640 19873 21649 19907
rect 21649 19873 21683 19907
rect 21683 19873 21692 19907
rect 21640 19864 21692 19873
rect 22100 19796 22152 19848
rect 21272 19660 21324 19712
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 20812 17824 20864 17876
rect 19984 17688 20036 17740
rect 21272 17731 21324 17740
rect 21272 17697 21281 17731
rect 21281 17697 21315 17731
rect 21315 17697 21324 17731
rect 21272 17688 21324 17697
rect 22744 17484 22796 17536
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 19984 14943 20036 14952
rect 19984 14909 19993 14943
rect 19993 14909 20027 14943
rect 20027 14909 20036 14943
rect 19984 14900 20036 14909
rect 20076 14764 20128 14816
rect 20260 14764 20312 14816
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 22744 14467 22796 14476
rect 22744 14433 22753 14467
rect 22753 14433 22787 14467
rect 22787 14433 22796 14467
rect 22744 14424 22796 14433
rect 23664 14220 23716 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 6644 12248 6696 12300
rect 20168 12291 20220 12300
rect 20168 12257 20177 12291
rect 20177 12257 20211 12291
rect 20211 12257 20220 12291
rect 20168 12248 20220 12257
rect 23664 12248 23716 12300
rect 24676 12248 24728 12300
rect 25412 12291 25464 12300
rect 25412 12257 25421 12291
rect 25421 12257 25455 12291
rect 25455 12257 25464 12291
rect 25412 12248 25464 12257
rect 23296 12112 23348 12164
rect 19432 12044 19484 12096
rect 19984 12087 20036 12096
rect 19984 12053 19993 12087
rect 19993 12053 20027 12087
rect 20027 12053 20036 12087
rect 19984 12044 20036 12053
rect 23388 12087 23440 12096
rect 23388 12053 23397 12087
rect 23397 12053 23431 12087
rect 23431 12053 23440 12087
rect 23388 12044 23440 12053
rect 25412 12044 25464 12096
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 22100 11840 22152 11892
rect 21548 11772 21600 11824
rect 20904 11636 20956 11688
rect 22376 11636 22428 11688
rect 22468 11568 22520 11620
rect 23664 11636 23716 11688
rect 25228 11636 25280 11688
rect 25412 11636 25464 11688
rect 27988 11636 28040 11688
rect 25596 11568 25648 11620
rect 23572 11500 23624 11552
rect 24124 11500 24176 11552
rect 24584 11500 24636 11552
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 20996 11228 21048 11280
rect 23388 11228 23440 11280
rect 23572 11203 23624 11212
rect 23572 11169 23581 11203
rect 23581 11169 23615 11203
rect 23615 11169 23624 11203
rect 23572 11160 23624 11169
rect 23664 11160 23716 11212
rect 25228 11203 25280 11212
rect 22652 11135 22704 11144
rect 22652 11101 22661 11135
rect 22661 11101 22695 11135
rect 22695 11101 22704 11135
rect 22652 11092 22704 11101
rect 23204 11092 23256 11144
rect 24768 11092 24820 11144
rect 21180 11067 21232 11076
rect 21180 11033 21189 11067
rect 21189 11033 21223 11067
rect 21223 11033 21232 11067
rect 21180 11024 21232 11033
rect 19708 10956 19760 11008
rect 20168 10956 20220 11008
rect 22284 10956 22336 11008
rect 23664 11024 23716 11076
rect 23204 10956 23256 11008
rect 24400 10956 24452 11008
rect 25228 11169 25237 11203
rect 25237 11169 25271 11203
rect 25271 11169 25280 11203
rect 25228 11160 25280 11169
rect 26240 11092 26292 11144
rect 25688 11024 25740 11076
rect 25780 11024 25832 11076
rect 26148 10956 26200 11008
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 22652 10752 22704 10804
rect 25596 10795 25648 10804
rect 25596 10761 25605 10795
rect 25605 10761 25639 10795
rect 25639 10761 25648 10795
rect 25596 10752 25648 10761
rect 30012 10752 30064 10804
rect 19064 10684 19116 10736
rect 19432 10548 19484 10600
rect 19708 10591 19760 10600
rect 19708 10557 19717 10591
rect 19717 10557 19751 10591
rect 19751 10557 19760 10591
rect 19708 10548 19760 10557
rect 19892 10548 19944 10600
rect 23572 10616 23624 10668
rect 27068 10616 27120 10668
rect 20812 10548 20864 10600
rect 22376 10548 22428 10600
rect 24400 10548 24452 10600
rect 24768 10548 24820 10600
rect 26240 10591 26292 10600
rect 22652 10480 22704 10532
rect 24676 10480 24728 10532
rect 26240 10557 26249 10591
rect 26249 10557 26283 10591
rect 26283 10557 26292 10591
rect 26240 10548 26292 10557
rect 19248 10412 19300 10464
rect 19340 10412 19392 10464
rect 20352 10412 20404 10464
rect 21272 10412 21324 10464
rect 22744 10412 22796 10464
rect 25964 10412 26016 10464
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 25780 10208 25832 10260
rect 19248 10140 19300 10192
rect 19432 10140 19484 10192
rect 19800 10072 19852 10124
rect 20352 10115 20404 10124
rect 20352 10081 20361 10115
rect 20361 10081 20395 10115
rect 20395 10081 20404 10115
rect 20352 10072 20404 10081
rect 18512 9868 18564 9920
rect 20904 10004 20956 10056
rect 20812 9979 20864 9988
rect 20812 9945 20821 9979
rect 20821 9945 20855 9979
rect 20855 9945 20864 9979
rect 20812 9936 20864 9945
rect 22928 10047 22980 10056
rect 22928 10013 22937 10047
rect 22937 10013 22971 10047
rect 22971 10013 22980 10047
rect 22928 10004 22980 10013
rect 23204 10047 23256 10056
rect 23204 10013 23213 10047
rect 23213 10013 23247 10047
rect 23247 10013 23256 10047
rect 23204 10004 23256 10013
rect 19248 9868 19300 9920
rect 20720 9868 20772 9920
rect 24676 10072 24728 10124
rect 24768 10072 24820 10124
rect 26148 10072 26200 10124
rect 26240 10072 26292 10124
rect 27160 10072 27212 10124
rect 27344 10115 27396 10124
rect 27344 10081 27353 10115
rect 27353 10081 27387 10115
rect 27387 10081 27396 10115
rect 27344 10072 27396 10081
rect 25228 10004 25280 10056
rect 25780 10004 25832 10056
rect 23756 9936 23808 9988
rect 24860 9868 24912 9920
rect 27160 9911 27212 9920
rect 27160 9877 27169 9911
rect 27169 9877 27203 9911
rect 27203 9877 27212 9911
rect 27160 9868 27212 9877
rect 31300 9868 31352 9920
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 17868 9528 17920 9580
rect 19800 9528 19852 9580
rect 20260 9528 20312 9580
rect 20628 9528 20680 9580
rect 22468 9596 22520 9648
rect 27804 9596 27856 9648
rect 24308 9528 24360 9580
rect 25228 9528 25280 9580
rect 27344 9528 27396 9580
rect 22100 9460 22152 9512
rect 22560 9503 22612 9512
rect 22560 9469 22569 9503
rect 22569 9469 22603 9503
rect 22603 9469 22612 9503
rect 22560 9460 22612 9469
rect 26516 9503 26568 9512
rect 26516 9469 26525 9503
rect 26525 9469 26559 9503
rect 26559 9469 26568 9503
rect 27988 9503 28040 9512
rect 26516 9460 26568 9469
rect 27988 9469 27997 9503
rect 27997 9469 28031 9503
rect 28031 9469 28040 9503
rect 27988 9460 28040 9469
rect 30380 9460 30432 9512
rect 19892 9392 19944 9444
rect 20168 9435 20220 9444
rect 20168 9401 20177 9435
rect 20177 9401 20211 9435
rect 20211 9401 20220 9435
rect 20168 9392 20220 9401
rect 22744 9392 22796 9444
rect 24952 9392 25004 9444
rect 25780 9392 25832 9444
rect 26240 9435 26292 9444
rect 26240 9401 26249 9435
rect 26249 9401 26283 9435
rect 26283 9401 26292 9435
rect 26240 9392 26292 9401
rect 28908 9392 28960 9444
rect 18696 9324 18748 9376
rect 21088 9324 21140 9376
rect 21732 9324 21784 9376
rect 22652 9324 22704 9376
rect 23848 9324 23900 9376
rect 25504 9324 25556 9376
rect 25596 9324 25648 9376
rect 28448 9367 28500 9376
rect 28448 9333 28457 9367
rect 28457 9333 28491 9367
rect 28491 9333 28500 9367
rect 28448 9324 28500 9333
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 19984 9052 20036 9104
rect 21548 9052 21600 9104
rect 22928 9120 22980 9172
rect 22376 9052 22428 9104
rect 24676 9120 24728 9172
rect 24952 9120 25004 9172
rect 24584 9052 24636 9104
rect 25504 9095 25556 9104
rect 25504 9061 25513 9095
rect 25513 9061 25547 9095
rect 25547 9061 25556 9095
rect 25504 9052 25556 9061
rect 26516 9052 26568 9104
rect 30472 9052 30524 9104
rect 17868 8984 17920 9036
rect 17224 8916 17276 8968
rect 20076 8984 20128 9036
rect 25136 8984 25188 9036
rect 27620 9027 27672 9036
rect 27620 8993 27629 9027
rect 27629 8993 27663 9027
rect 27663 8993 27672 9027
rect 27620 8984 27672 8993
rect 28908 9027 28960 9036
rect 19432 8916 19484 8968
rect 18328 8780 18380 8832
rect 21732 8916 21784 8968
rect 22468 8959 22520 8968
rect 22468 8925 22477 8959
rect 22477 8925 22511 8959
rect 22511 8925 22520 8959
rect 22468 8916 22520 8925
rect 22744 8959 22796 8968
rect 22744 8925 22753 8959
rect 22753 8925 22787 8959
rect 22787 8925 22796 8959
rect 22744 8916 22796 8925
rect 28908 8993 28917 9027
rect 28917 8993 28951 9027
rect 28951 8993 28960 9027
rect 28908 8984 28960 8993
rect 20628 8780 20680 8832
rect 20904 8780 20956 8832
rect 27712 8848 27764 8900
rect 30196 8916 30248 8968
rect 24216 8823 24268 8832
rect 24216 8789 24225 8823
rect 24225 8789 24259 8823
rect 24259 8789 24268 8823
rect 24216 8780 24268 8789
rect 26608 8780 26660 8832
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 17316 8576 17368 8628
rect 20076 8576 20128 8628
rect 21272 8576 21324 8628
rect 22192 8576 22244 8628
rect 24860 8576 24912 8628
rect 25780 8576 25832 8628
rect 26516 8619 26568 8628
rect 26516 8585 26525 8619
rect 26525 8585 26559 8619
rect 26559 8585 26568 8619
rect 26516 8576 26568 8585
rect 17960 8440 18012 8492
rect 19432 8415 19484 8424
rect 19432 8381 19441 8415
rect 19441 8381 19475 8415
rect 19475 8381 19484 8415
rect 22928 8440 22980 8492
rect 25596 8508 25648 8560
rect 19432 8372 19484 8381
rect 22560 8372 22612 8424
rect 25228 8415 25280 8424
rect 25228 8381 25237 8415
rect 25237 8381 25271 8415
rect 25271 8381 25280 8415
rect 25228 8372 25280 8381
rect 18696 8304 18748 8356
rect 20904 8304 20956 8356
rect 17684 8279 17736 8288
rect 17684 8245 17693 8279
rect 17693 8245 17727 8279
rect 17727 8245 17736 8279
rect 17684 8236 17736 8245
rect 18788 8236 18840 8288
rect 23572 8304 23624 8356
rect 25044 8304 25096 8356
rect 25320 8236 25372 8288
rect 27344 8372 27396 8424
rect 26792 8304 26844 8356
rect 29184 8372 29236 8424
rect 30380 8372 30432 8424
rect 31484 8372 31536 8424
rect 25780 8236 25832 8288
rect 29552 8279 29604 8288
rect 29552 8245 29561 8279
rect 29561 8245 29595 8279
rect 29595 8245 29604 8279
rect 29552 8236 29604 8245
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 14924 7760 14976 7812
rect 16212 7896 16264 7948
rect 17224 7896 17276 7948
rect 17684 7964 17736 8016
rect 20168 8032 20220 8084
rect 20260 8032 20312 8084
rect 23480 8032 23532 8084
rect 23572 8032 23624 8084
rect 26240 8032 26292 8084
rect 22928 7964 22980 8016
rect 25780 7964 25832 8016
rect 30288 8032 30340 8084
rect 29552 7964 29604 8016
rect 18696 7896 18748 7948
rect 19432 7896 19484 7948
rect 19892 7896 19944 7948
rect 27344 7896 27396 7948
rect 29276 7896 29328 7948
rect 31300 7939 31352 7948
rect 19340 7828 19392 7880
rect 22560 7871 22612 7880
rect 22560 7837 22569 7871
rect 22569 7837 22603 7871
rect 22603 7837 22612 7871
rect 22560 7828 22612 7837
rect 22836 7871 22888 7880
rect 22836 7837 22845 7871
rect 22845 7837 22879 7871
rect 22879 7837 22888 7871
rect 22836 7828 22888 7837
rect 23480 7828 23532 7880
rect 15108 7692 15160 7744
rect 16672 7735 16724 7744
rect 16672 7701 16681 7735
rect 16681 7701 16715 7735
rect 16715 7701 16724 7735
rect 16672 7692 16724 7701
rect 16764 7692 16816 7744
rect 20996 7692 21048 7744
rect 22376 7692 22428 7744
rect 24952 7692 25004 7744
rect 25136 7828 25188 7880
rect 25504 7871 25556 7880
rect 25504 7837 25513 7871
rect 25513 7837 25547 7871
rect 25547 7837 25556 7871
rect 25504 7828 25556 7837
rect 25596 7828 25648 7880
rect 28908 7828 28960 7880
rect 31300 7905 31309 7939
rect 31309 7905 31343 7939
rect 31343 7905 31352 7939
rect 31300 7896 31352 7905
rect 26608 7692 26660 7744
rect 26792 7692 26844 7744
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 16764 7488 16816 7540
rect 16580 7420 16632 7472
rect 15200 7352 15252 7404
rect 22836 7488 22888 7540
rect 24124 7488 24176 7540
rect 24952 7531 25004 7540
rect 24952 7497 24961 7531
rect 24961 7497 24995 7531
rect 24995 7497 25004 7531
rect 24952 7488 25004 7497
rect 25320 7488 25372 7540
rect 28632 7488 28684 7540
rect 29184 7488 29236 7540
rect 30196 7463 30248 7472
rect 30196 7429 30205 7463
rect 30205 7429 30239 7463
rect 30239 7429 30248 7463
rect 30196 7420 30248 7429
rect 19432 7352 19484 7404
rect 20536 7352 20588 7404
rect 23664 7352 23716 7404
rect 24216 7395 24268 7404
rect 24216 7361 24225 7395
rect 24225 7361 24259 7395
rect 24259 7361 24268 7395
rect 24216 7352 24268 7361
rect 24492 7395 24544 7404
rect 24492 7361 24501 7395
rect 24501 7361 24535 7395
rect 24535 7361 24544 7395
rect 24492 7352 24544 7361
rect 25412 7352 25464 7404
rect 26700 7395 26752 7404
rect 26700 7361 26709 7395
rect 26709 7361 26743 7395
rect 26743 7361 26752 7395
rect 26700 7352 26752 7361
rect 27712 7352 27764 7404
rect 28172 7352 28224 7404
rect 29276 7352 29328 7404
rect 29552 7352 29604 7404
rect 14924 7327 14976 7336
rect 14924 7293 14933 7327
rect 14933 7293 14967 7327
rect 14967 7293 14976 7327
rect 14924 7284 14976 7293
rect 15016 7284 15068 7336
rect 16212 7327 16264 7336
rect 16212 7293 16221 7327
rect 16221 7293 16255 7327
rect 16255 7293 16264 7327
rect 16212 7284 16264 7293
rect 19892 7327 19944 7336
rect 19892 7293 19901 7327
rect 19901 7293 19935 7327
rect 19935 7293 19944 7327
rect 19892 7284 19944 7293
rect 30012 7327 30064 7336
rect 17868 7216 17920 7268
rect 20444 7216 20496 7268
rect 22652 7216 22704 7268
rect 17500 7148 17552 7200
rect 19984 7148 20036 7200
rect 21640 7191 21692 7200
rect 21640 7157 21649 7191
rect 21649 7157 21683 7191
rect 21683 7157 21692 7191
rect 21640 7148 21692 7157
rect 25964 7216 26016 7268
rect 30012 7293 30021 7327
rect 30021 7293 30055 7327
rect 30055 7293 30064 7327
rect 30012 7284 30064 7293
rect 30840 7327 30892 7336
rect 30840 7293 30849 7327
rect 30849 7293 30883 7327
rect 30883 7293 30892 7327
rect 30840 7284 30892 7293
rect 31484 7327 31536 7336
rect 31484 7293 31493 7327
rect 31493 7293 31527 7327
rect 31527 7293 31536 7327
rect 31484 7284 31536 7293
rect 28172 7216 28224 7268
rect 29828 7216 29880 7268
rect 27160 7148 27212 7200
rect 28724 7148 28776 7200
rect 30380 7148 30432 7200
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 15108 6944 15160 6996
rect 20168 6987 20220 6996
rect 16028 6876 16080 6928
rect 14648 6808 14700 6860
rect 15108 6851 15160 6860
rect 15108 6817 15117 6851
rect 15117 6817 15151 6851
rect 15151 6817 15160 6851
rect 15108 6808 15160 6817
rect 20168 6953 20177 6987
rect 20177 6953 20211 6987
rect 20211 6953 20220 6987
rect 20168 6944 20220 6953
rect 20260 6876 20312 6928
rect 21640 6919 21692 6928
rect 21640 6885 21649 6919
rect 21649 6885 21683 6919
rect 21683 6885 21692 6919
rect 21640 6876 21692 6885
rect 23296 6876 23348 6928
rect 24124 6944 24176 6996
rect 25320 6876 25372 6928
rect 25688 6876 25740 6928
rect 26700 6876 26752 6928
rect 16764 6808 16816 6860
rect 22560 6808 22612 6860
rect 24400 6808 24452 6860
rect 27804 6876 27856 6928
rect 30012 6876 30064 6928
rect 27436 6851 27488 6860
rect 27436 6817 27445 6851
rect 27445 6817 27479 6851
rect 27479 6817 27488 6851
rect 27436 6808 27488 6817
rect 30472 6808 30524 6860
rect 31300 6876 31352 6928
rect 15384 6783 15436 6792
rect 15384 6749 15393 6783
rect 15393 6749 15427 6783
rect 15427 6749 15436 6783
rect 15384 6740 15436 6749
rect 16580 6740 16632 6792
rect 22468 6740 22520 6792
rect 23848 6783 23900 6792
rect 23848 6749 23857 6783
rect 23857 6749 23891 6783
rect 23891 6749 23900 6783
rect 23848 6740 23900 6749
rect 24952 6740 25004 6792
rect 20628 6672 20680 6724
rect 22744 6672 22796 6724
rect 27252 6672 27304 6724
rect 16856 6647 16908 6656
rect 16856 6613 16865 6647
rect 16865 6613 16899 6647
rect 16899 6613 16908 6647
rect 16856 6604 16908 6613
rect 16948 6604 17000 6656
rect 21180 6604 21232 6656
rect 22836 6604 22888 6656
rect 26148 6604 26200 6656
rect 28816 6604 28868 6656
rect 29368 6604 29420 6656
rect 30840 6604 30892 6656
rect 31668 6604 31720 6656
rect 32404 6647 32456 6656
rect 32404 6613 32413 6647
rect 32413 6613 32447 6647
rect 32447 6613 32456 6647
rect 32404 6604 32456 6613
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 15384 6400 15436 6452
rect 16856 6400 16908 6452
rect 16028 6264 16080 6316
rect 16948 6332 17000 6384
rect 19432 6375 19484 6384
rect 19432 6341 19441 6375
rect 19441 6341 19475 6375
rect 19475 6341 19484 6375
rect 19432 6332 19484 6341
rect 22192 6400 22244 6452
rect 24308 6443 24360 6452
rect 16580 6264 16632 6316
rect 17960 6307 18012 6316
rect 15200 6060 15252 6112
rect 16672 6060 16724 6112
rect 17960 6273 17969 6307
rect 17969 6273 18003 6307
rect 18003 6273 18012 6307
rect 17960 6264 18012 6273
rect 19156 6264 19208 6316
rect 19892 6239 19944 6248
rect 19892 6205 19901 6239
rect 19901 6205 19935 6239
rect 19935 6205 19944 6239
rect 19892 6196 19944 6205
rect 21456 6196 21508 6248
rect 22192 6196 22244 6248
rect 22376 6264 22428 6316
rect 24308 6409 24317 6443
rect 24317 6409 24351 6443
rect 24351 6409 24360 6443
rect 24308 6400 24360 6409
rect 24860 6400 24912 6452
rect 26792 6400 26844 6452
rect 27252 6400 27304 6452
rect 29828 6400 29880 6452
rect 30288 6400 30340 6452
rect 30472 6332 30524 6384
rect 22560 6239 22612 6248
rect 19340 6060 19392 6112
rect 20168 6171 20220 6180
rect 20168 6137 20177 6171
rect 20177 6137 20211 6171
rect 20211 6137 20220 6171
rect 20168 6128 20220 6137
rect 21456 6060 21508 6112
rect 21824 6128 21876 6180
rect 22284 6128 22336 6180
rect 22100 6060 22152 6112
rect 22560 6205 22569 6239
rect 22569 6205 22603 6239
rect 22603 6205 22612 6239
rect 22560 6196 22612 6205
rect 24860 6196 24912 6248
rect 26516 6239 26568 6248
rect 26516 6205 26525 6239
rect 26525 6205 26559 6239
rect 26559 6205 26568 6239
rect 26516 6196 26568 6205
rect 27436 6196 27488 6248
rect 29368 6196 29420 6248
rect 30288 6196 30340 6248
rect 24768 6103 24820 6112
rect 24768 6069 24777 6103
rect 24777 6069 24811 6103
rect 24811 6069 24820 6103
rect 24768 6060 24820 6069
rect 26148 6128 26200 6180
rect 26976 6128 27028 6180
rect 28172 6060 28224 6112
rect 31668 6128 31720 6180
rect 31944 6103 31996 6112
rect 31944 6069 31953 6103
rect 31953 6069 31987 6103
rect 31987 6069 31996 6103
rect 31944 6060 31996 6069
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 17316 5899 17368 5908
rect 17316 5865 17325 5899
rect 17325 5865 17359 5899
rect 17359 5865 17368 5899
rect 17316 5856 17368 5865
rect 21548 5856 21600 5908
rect 24124 5856 24176 5908
rect 25412 5856 25464 5908
rect 26976 5899 27028 5908
rect 26976 5865 26985 5899
rect 26985 5865 27019 5899
rect 27019 5865 27028 5899
rect 26976 5856 27028 5865
rect 22836 5788 22888 5840
rect 23756 5788 23808 5840
rect 24860 5788 24912 5840
rect 30380 5856 30432 5908
rect 28448 5788 28500 5840
rect 28816 5788 28868 5840
rect 15016 5720 15068 5772
rect 16856 5763 16908 5772
rect 16856 5729 16865 5763
rect 16865 5729 16899 5763
rect 16899 5729 16908 5763
rect 16856 5720 16908 5729
rect 19340 5720 19392 5772
rect 22468 5763 22520 5772
rect 22468 5729 22477 5763
rect 22477 5729 22511 5763
rect 22511 5729 22520 5763
rect 22468 5720 22520 5729
rect 24400 5720 24452 5772
rect 25228 5763 25280 5772
rect 25228 5729 25237 5763
rect 25237 5729 25271 5763
rect 25271 5729 25280 5763
rect 25228 5720 25280 5729
rect 29276 5720 29328 5772
rect 18788 5695 18840 5704
rect 18788 5661 18797 5695
rect 18797 5661 18831 5695
rect 18831 5661 18840 5695
rect 18788 5652 18840 5661
rect 22284 5652 22336 5704
rect 28172 5652 28224 5704
rect 28356 5652 28408 5704
rect 30012 5652 30064 5704
rect 31392 5788 31444 5840
rect 31668 5788 31720 5840
rect 31300 5720 31352 5772
rect 32404 5652 32456 5704
rect 15108 5559 15160 5568
rect 15108 5525 15117 5559
rect 15117 5525 15151 5559
rect 15151 5525 15160 5559
rect 15108 5516 15160 5525
rect 22836 5516 22888 5568
rect 24124 5516 24176 5568
rect 27436 5559 27488 5568
rect 27436 5525 27445 5559
rect 27445 5525 27479 5559
rect 27479 5525 27488 5559
rect 27436 5516 27488 5525
rect 29368 5584 29420 5636
rect 30288 5584 30340 5636
rect 28172 5516 28224 5568
rect 28264 5516 28316 5568
rect 30472 5559 30524 5568
rect 30472 5525 30481 5559
rect 30481 5525 30515 5559
rect 30515 5525 30524 5559
rect 31300 5559 31352 5568
rect 30472 5516 30524 5525
rect 31300 5525 31309 5559
rect 31309 5525 31343 5559
rect 31343 5525 31352 5559
rect 31300 5516 31352 5525
rect 31760 5559 31812 5568
rect 31760 5525 31769 5559
rect 31769 5525 31803 5559
rect 31803 5525 31812 5559
rect 31760 5516 31812 5525
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 18788 5312 18840 5364
rect 24860 5355 24912 5364
rect 24860 5321 24869 5355
rect 24869 5321 24903 5355
rect 24903 5321 24912 5355
rect 24860 5312 24912 5321
rect 24952 5244 25004 5296
rect 16488 5176 16540 5228
rect 19432 5219 19484 5228
rect 19432 5185 19441 5219
rect 19441 5185 19475 5219
rect 19475 5185 19484 5219
rect 19432 5176 19484 5185
rect 21180 5176 21232 5228
rect 22560 5176 22612 5228
rect 24768 5176 24820 5228
rect 14648 5151 14700 5160
rect 14648 5117 14657 5151
rect 14657 5117 14691 5151
rect 14691 5117 14700 5151
rect 14648 5108 14700 5117
rect 14924 5083 14976 5092
rect 14924 5049 14933 5083
rect 14933 5049 14967 5083
rect 14967 5049 14976 5083
rect 14924 5040 14976 5049
rect 17868 5040 17920 5092
rect 19064 5040 19116 5092
rect 20076 5040 20128 5092
rect 15108 4972 15160 5024
rect 17592 4972 17644 5024
rect 22376 4972 22428 5024
rect 24032 5108 24084 5160
rect 25872 5176 25924 5228
rect 28264 5244 28316 5296
rect 30380 5244 30432 5296
rect 26700 5176 26752 5228
rect 26332 5083 26384 5092
rect 26332 5049 26341 5083
rect 26341 5049 26375 5083
rect 26375 5049 26384 5083
rect 26332 5040 26384 5049
rect 31944 5176 31996 5228
rect 29552 5151 29604 5160
rect 29552 5117 29561 5151
rect 29561 5117 29595 5151
rect 29595 5117 29604 5151
rect 29552 5108 29604 5117
rect 30012 5108 30064 5160
rect 30656 5108 30708 5160
rect 31300 5108 31352 5160
rect 27988 5040 28040 5092
rect 29276 5083 29328 5092
rect 29276 5049 29285 5083
rect 29285 5049 29319 5083
rect 29319 5049 29328 5083
rect 29276 5040 29328 5049
rect 27896 4972 27948 5024
rect 28908 4972 28960 5024
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 14924 4768 14976 4820
rect 17868 4768 17920 4820
rect 16120 4700 16172 4752
rect 18328 4700 18380 4752
rect 22836 4743 22888 4752
rect 16856 4675 16908 4684
rect 16856 4641 16865 4675
rect 16865 4641 16899 4675
rect 16899 4641 16908 4675
rect 17316 4675 17368 4684
rect 16856 4632 16908 4641
rect 17316 4641 17325 4675
rect 17325 4641 17359 4675
rect 17359 4641 17368 4675
rect 17316 4632 17368 4641
rect 16580 4607 16632 4616
rect 16580 4573 16589 4607
rect 16589 4573 16623 4607
rect 16623 4573 16632 4607
rect 16580 4564 16632 4573
rect 17684 4564 17736 4616
rect 22836 4709 22845 4743
rect 22845 4709 22879 4743
rect 22879 4709 22888 4743
rect 22836 4700 22888 4709
rect 25872 4700 25924 4752
rect 26240 4700 26292 4752
rect 29276 4768 29328 4820
rect 22560 4675 22612 4684
rect 20720 4564 20772 4616
rect 22560 4641 22569 4675
rect 22569 4641 22603 4675
rect 22603 4641 22612 4675
rect 22560 4632 22612 4641
rect 27804 4632 27856 4684
rect 20628 4496 20680 4548
rect 19892 4428 19944 4480
rect 19984 4428 20036 4480
rect 20444 4428 20496 4480
rect 26700 4564 26752 4616
rect 26792 4564 26844 4616
rect 28724 4700 28776 4752
rect 29184 4675 29236 4684
rect 29184 4641 29193 4675
rect 29193 4641 29227 4675
rect 29227 4641 29236 4675
rect 29184 4632 29236 4641
rect 30656 4675 30708 4684
rect 30656 4641 30665 4675
rect 30665 4641 30699 4675
rect 30699 4641 30708 4675
rect 30656 4632 30708 4641
rect 28264 4564 28316 4616
rect 26608 4428 26660 4480
rect 26700 4428 26752 4480
rect 28356 4428 28408 4480
rect 30472 4471 30524 4480
rect 30472 4437 30481 4471
rect 30481 4437 30515 4471
rect 30515 4437 30524 4471
rect 30472 4428 30524 4437
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 16120 4224 16172 4276
rect 16580 4224 16632 4276
rect 17776 4224 17828 4276
rect 19984 4224 20036 4276
rect 22928 4224 22980 4276
rect 27436 4224 27488 4276
rect 27804 4267 27856 4276
rect 27804 4233 27813 4267
rect 27813 4233 27847 4267
rect 27847 4233 27856 4267
rect 27804 4224 27856 4233
rect 17316 4088 17368 4140
rect 18512 4088 18564 4140
rect 18604 4088 18656 4140
rect 23112 4156 23164 4208
rect 22284 4088 22336 4140
rect 24860 4088 24912 4140
rect 30472 4156 30524 4208
rect 16120 4020 16172 4072
rect 16396 4063 16448 4072
rect 16396 4029 16405 4063
rect 16405 4029 16439 4063
rect 16439 4029 16448 4063
rect 16396 4020 16448 4029
rect 19432 4020 19484 4072
rect 27620 4088 27672 4140
rect 27896 4088 27948 4140
rect 17960 3995 18012 4004
rect 17684 3884 17736 3936
rect 17960 3961 17969 3995
rect 17969 3961 18003 3995
rect 18003 3961 18012 3995
rect 17960 3952 18012 3961
rect 19248 3952 19300 4004
rect 20444 3952 20496 4004
rect 22836 3952 22888 4004
rect 23664 3952 23716 4004
rect 24216 3952 24268 4004
rect 25228 3952 25280 4004
rect 21456 3884 21508 3936
rect 22468 3884 22520 3936
rect 22652 3884 22704 3936
rect 27896 3952 27948 4004
rect 28172 4020 28224 4072
rect 29368 4020 29420 4072
rect 30656 4088 30708 4140
rect 28264 3952 28316 4004
rect 26700 3927 26752 3936
rect 26700 3893 26709 3927
rect 26709 3893 26743 3927
rect 26743 3893 26752 3927
rect 26700 3884 26752 3893
rect 28632 3884 28684 3936
rect 29000 3884 29052 3936
rect 29644 3884 29696 3936
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 15752 3544 15804 3596
rect 16580 3612 16632 3664
rect 17592 3655 17644 3664
rect 17592 3621 17601 3655
rect 17601 3621 17635 3655
rect 17635 3621 17644 3655
rect 17592 3612 17644 3621
rect 18604 3612 18656 3664
rect 22376 3612 22428 3664
rect 24216 3680 24268 3732
rect 24584 3680 24636 3732
rect 27068 3680 27120 3732
rect 27620 3680 27672 3732
rect 29000 3612 29052 3664
rect 16120 3544 16172 3596
rect 17316 3587 17368 3596
rect 17316 3553 17325 3587
rect 17325 3553 17359 3587
rect 17359 3553 17368 3587
rect 17316 3544 17368 3553
rect 22192 3544 22244 3596
rect 22560 3587 22612 3596
rect 22560 3553 22569 3587
rect 22569 3553 22603 3587
rect 22603 3553 22612 3587
rect 22560 3544 22612 3553
rect 24860 3544 24912 3596
rect 25228 3587 25280 3596
rect 25228 3553 25237 3587
rect 25237 3553 25271 3587
rect 25271 3553 25280 3587
rect 25228 3544 25280 3553
rect 27252 3544 27304 3596
rect 27344 3544 27396 3596
rect 28172 3544 28224 3596
rect 28540 3544 28592 3596
rect 28908 3587 28960 3596
rect 28908 3553 28917 3587
rect 28917 3553 28951 3587
rect 28951 3553 28960 3587
rect 28908 3544 28960 3553
rect 29552 3587 29604 3596
rect 29552 3553 29561 3587
rect 29561 3553 29595 3587
rect 29595 3553 29604 3587
rect 29552 3544 29604 3553
rect 31392 3544 31444 3596
rect 19432 3476 19484 3528
rect 18052 3340 18104 3392
rect 20352 3383 20404 3392
rect 20352 3349 20361 3383
rect 20361 3349 20395 3383
rect 20395 3349 20404 3383
rect 20352 3340 20404 3349
rect 26792 3476 26844 3528
rect 27896 3476 27948 3528
rect 27988 3408 28040 3460
rect 28356 3476 28408 3528
rect 31760 3408 31812 3460
rect 22836 3340 22888 3392
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 17776 3136 17828 3188
rect 17960 3136 18012 3188
rect 19432 3179 19484 3188
rect 19432 3145 19441 3179
rect 19441 3145 19475 3179
rect 19475 3145 19484 3179
rect 19432 3136 19484 3145
rect 20076 3136 20128 3188
rect 21180 3136 21232 3188
rect 26332 3136 26384 3188
rect 26608 3179 26660 3188
rect 26608 3145 26617 3179
rect 26617 3145 26651 3179
rect 26651 3145 26660 3179
rect 26608 3136 26660 3145
rect 26884 3136 26936 3188
rect 26976 3136 27028 3188
rect 29184 3136 29236 3188
rect 17500 3068 17552 3120
rect 15108 2932 15160 2984
rect 18052 2975 18104 2984
rect 18052 2941 18061 2975
rect 18061 2941 18095 2975
rect 18095 2941 18104 2975
rect 18052 2932 18104 2941
rect 16488 2864 16540 2916
rect 18696 2932 18748 2984
rect 19156 2975 19208 2984
rect 19156 2941 19165 2975
rect 19165 2941 19199 2975
rect 19199 2941 19208 2975
rect 19156 2932 19208 2941
rect 26240 3068 26292 3120
rect 27068 3068 27120 3120
rect 20628 3000 20680 3052
rect 22192 3000 22244 3052
rect 22468 3000 22520 3052
rect 24676 2932 24728 2984
rect 24584 2864 24636 2916
rect 11152 2839 11204 2848
rect 11152 2805 11161 2839
rect 11161 2805 11195 2839
rect 11195 2805 11204 2839
rect 11152 2796 11204 2805
rect 16396 2796 16448 2848
rect 25780 2932 25832 2984
rect 29644 3000 29696 3052
rect 26700 2975 26752 2984
rect 26700 2941 26709 2975
rect 26709 2941 26743 2975
rect 26743 2941 26752 2975
rect 26700 2932 26752 2941
rect 28356 2932 28408 2984
rect 29552 2932 29604 2984
rect 28264 2864 28316 2916
rect 28724 2864 28776 2916
rect 25044 2796 25096 2848
rect 28448 2839 28500 2848
rect 28448 2805 28457 2839
rect 28457 2805 28491 2839
rect 28491 2805 28500 2839
rect 28448 2796 28500 2805
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 20720 2592 20772 2644
rect 22928 2635 22980 2644
rect 22928 2601 22937 2635
rect 22937 2601 22971 2635
rect 22971 2601 22980 2635
rect 22928 2592 22980 2601
rect 23112 2592 23164 2644
rect 25780 2592 25832 2644
rect 11152 2524 11204 2576
rect 15752 2567 15804 2576
rect 15752 2533 15761 2567
rect 15761 2533 15795 2567
rect 15795 2533 15804 2567
rect 15752 2524 15804 2533
rect 18696 2567 18748 2576
rect 18696 2533 18705 2567
rect 18705 2533 18739 2567
rect 18739 2533 18748 2567
rect 18696 2524 18748 2533
rect 21088 2524 21140 2576
rect 21456 2524 21508 2576
rect 25044 2524 25096 2576
rect 26608 2592 26660 2644
rect 26884 2592 26936 2644
rect 20352 2456 20404 2508
rect 22284 2456 22336 2508
rect 25228 2456 25280 2508
rect 26976 2524 27028 2576
rect 28264 2592 28316 2644
rect 20260 2431 20312 2440
rect 20260 2397 20269 2431
rect 20269 2397 20303 2431
rect 20303 2397 20312 2431
rect 20260 2388 20312 2397
rect 26792 2456 26844 2508
rect 28356 2456 28408 2508
rect 2228 2363 2280 2372
rect 2228 2329 2237 2363
rect 2237 2329 2271 2363
rect 2271 2329 2280 2363
rect 2228 2320 2280 2329
rect 11060 2363 11112 2372
rect 11060 2329 11069 2363
rect 11069 2329 11103 2363
rect 11103 2329 11112 2363
rect 11060 2320 11112 2329
rect 15568 2363 15620 2372
rect 15568 2329 15577 2363
rect 15577 2329 15611 2363
rect 15611 2329 15620 2363
rect 15568 2320 15620 2329
rect 19984 2320 20036 2372
rect 28172 2388 28224 2440
rect 27068 2320 27120 2372
rect 28908 2363 28960 2372
rect 28908 2329 28917 2363
rect 28917 2329 28951 2363
rect 28951 2329 28960 2363
rect 28908 2320 28960 2329
rect 33324 2320 33376 2372
rect 37740 2363 37792 2372
rect 37740 2329 37749 2363
rect 37749 2329 37783 2363
rect 37783 2329 37792 2363
rect 37740 2320 37792 2329
rect 22100 2252 22152 2304
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
rect 24400 960 24452 1012
rect 28724 960 28776 1012
<< metal2 >>
rect 19982 39200 20038 40000
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 19996 36718 20024 39200
rect 20812 37324 20864 37330
rect 20812 37266 20864 37272
rect 20444 37256 20496 37262
rect 20444 37198 20496 37204
rect 20456 36922 20484 37198
rect 20444 36916 20496 36922
rect 20444 36858 20496 36864
rect 19984 36712 20036 36718
rect 19984 36654 20036 36660
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 19984 21548 20036 21554
rect 19984 21490 20036 21496
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 19076 21010 19104 21422
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19996 21010 20024 21490
rect 20824 21418 20852 37266
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 20812 21412 20864 21418
rect 20812 21354 20864 21360
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 20364 21010 20392 21286
rect 20824 21146 20852 21354
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 19064 21004 19116 21010
rect 19064 20946 19116 20952
rect 19984 21004 20036 21010
rect 19984 20946 20036 20952
rect 20352 21004 20404 21010
rect 20352 20946 20404 20952
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 19996 20466 20024 20946
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 19996 17746 20024 20402
rect 20824 20330 20852 21082
rect 20904 20800 20956 20806
rect 20904 20742 20956 20748
rect 20916 20466 20944 20742
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 20904 20460 20956 20466
rect 20904 20402 20956 20408
rect 20812 20324 20864 20330
rect 20812 20266 20864 20272
rect 20824 19990 20852 20266
rect 21640 20256 21692 20262
rect 21640 20198 21692 20204
rect 20812 19984 20864 19990
rect 20812 19926 20864 19932
rect 20824 17882 20852 19926
rect 21652 19922 21680 20198
rect 21640 19916 21692 19922
rect 21640 19858 21692 19864
rect 22100 19848 22152 19854
rect 22100 19790 22152 19796
rect 21272 19712 21324 19718
rect 21272 19654 21324 19660
rect 20812 17876 20864 17882
rect 20812 17818 20864 17824
rect 21284 17746 21312 19654
rect 19984 17740 20036 17746
rect 19984 17682 20036 17688
rect 21272 17740 21324 17746
rect 21272 17682 21324 17688
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19996 16574 20024 17682
rect 19996 16546 20116 16574
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 6644 12300 6696 12306
rect 6644 12242 6696 12248
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 2228 2372 2280 2378
rect 2228 2314 2280 2320
rect 2240 800 2268 2314
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 6656 800 6684 12242
rect 19996 12102 20024 14894
rect 20088 14822 20116 16546
rect 20076 14816 20128 14822
rect 20076 14758 20128 14764
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 20168 12300 20220 12306
rect 20168 12242 20220 12248
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 19064 10736 19116 10742
rect 19064 10678 19116 10684
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 17880 9042 17908 9522
rect 17868 9036 17920 9042
rect 17868 8978 17920 8984
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17236 7954 17264 8910
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 14924 7812 14976 7818
rect 14924 7754 14976 7760
rect 14936 7342 14964 7754
rect 15108 7744 15160 7750
rect 15108 7686 15160 7692
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14660 5166 14688 6802
rect 15028 5778 15056 7278
rect 15120 7002 15148 7686
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 15120 6866 15148 6938
rect 15108 6860 15160 6866
rect 15108 6802 15160 6808
rect 15212 6118 15240 7346
rect 16224 7342 16252 7890
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16580 7472 16632 7478
rect 16580 7414 16632 7420
rect 16212 7336 16264 7342
rect 16212 7278 16264 7284
rect 16028 6928 16080 6934
rect 16028 6870 16080 6876
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 15396 6458 15424 6734
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 16040 6322 16068 6870
rect 16592 6798 16620 7414
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 16592 6322 16620 6734
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 16684 6118 16712 7686
rect 16776 7546 16804 7686
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16764 6860 16816 6866
rect 16764 6802 16816 6808
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 15016 5772 15068 5778
rect 16776 5760 16804 6802
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16868 6458 16896 6598
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16960 6390 16988 6598
rect 16948 6384 17000 6390
rect 16948 6326 17000 6332
rect 17328 5914 17356 8570
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17696 8022 17724 8230
rect 17684 8016 17736 8022
rect 17684 7958 17736 7964
rect 17880 7274 17908 8978
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17868 7268 17920 7274
rect 17868 7210 17920 7216
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 16856 5772 16908 5778
rect 16776 5732 16856 5760
rect 15016 5714 15068 5720
rect 16856 5714 16908 5720
rect 15108 5568 15160 5574
rect 15108 5510 15160 5516
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14924 5092 14976 5098
rect 14924 5034 14976 5040
rect 14936 4826 14964 5034
rect 15120 5030 15148 5510
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 15108 5024 15160 5030
rect 15108 4966 15160 4972
rect 14924 4820 14976 4826
rect 14924 4762 14976 4768
rect 15120 2990 15148 4966
rect 16120 4752 16172 4758
rect 16120 4694 16172 4700
rect 16132 4282 16160 4694
rect 16120 4276 16172 4282
rect 16120 4218 16172 4224
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16132 3602 16160 4014
rect 15752 3596 15804 3602
rect 15752 3538 15804 3544
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 15108 2984 15160 2990
rect 15108 2926 15160 2932
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 11164 2582 11192 2790
rect 15764 2582 15792 3538
rect 16408 2854 16436 4014
rect 16500 2922 16528 5170
rect 16868 4690 16896 5714
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16592 4282 16620 4558
rect 16580 4276 16632 4282
rect 16580 4218 16632 4224
rect 16592 3670 16620 4218
rect 17328 4146 17356 4626
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 16580 3664 16632 3670
rect 16580 3606 16632 3612
rect 17328 3602 17356 4082
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 17512 3126 17540 7142
rect 17972 6322 18000 8434
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 17868 5092 17920 5098
rect 17868 5034 17920 5040
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 17604 3670 17632 4966
rect 17880 4826 17908 5034
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 18340 4758 18368 8774
rect 18328 4752 18380 4758
rect 18328 4694 18380 4700
rect 17684 4616 17736 4622
rect 17684 4558 17736 4564
rect 17696 3942 17724 4558
rect 17776 4276 17828 4282
rect 17776 4218 17828 4224
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17592 3664 17644 3670
rect 17592 3606 17644 3612
rect 17788 3194 17816 4218
rect 18524 4146 18552 9862
rect 18696 9376 18748 9382
rect 18696 9318 18748 9324
rect 18708 8362 18736 9318
rect 18696 8356 18748 8362
rect 18696 8298 18748 8304
rect 18788 8288 18840 8294
rect 18788 8230 18840 8236
rect 18800 8106 18828 8230
rect 18708 8078 18828 8106
rect 18708 7954 18736 8078
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18800 5370 18828 5646
rect 18788 5364 18840 5370
rect 18788 5306 18840 5312
rect 19076 5098 19104 10678
rect 19444 10606 19472 12038
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 20180 11014 20208 12242
rect 19708 11008 19760 11014
rect 19708 10950 19760 10956
rect 20168 11008 20220 11014
rect 20168 10950 20220 10956
rect 19720 10606 19748 10950
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19892 10600 19944 10606
rect 19892 10542 19944 10548
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19260 10198 19288 10406
rect 19248 10192 19300 10198
rect 19248 10134 19300 10140
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 19064 5092 19116 5098
rect 19064 5034 19116 5040
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 17960 4004 18012 4010
rect 17960 3946 18012 3952
rect 17972 3194 18000 3946
rect 18616 3670 18644 4082
rect 18604 3664 18656 3670
rect 18604 3606 18656 3612
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 17500 3120 17552 3126
rect 17500 3062 17552 3068
rect 18064 2990 18092 3334
rect 19168 2990 19196 6258
rect 19260 4010 19288 9862
rect 19352 7886 19380 10406
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 19432 10192 19484 10198
rect 19432 10134 19484 10140
rect 19444 8974 19472 10134
rect 19800 10124 19852 10130
rect 19800 10066 19852 10072
rect 19812 9586 19840 10066
rect 19800 9580 19852 9586
rect 19800 9522 19852 9528
rect 19904 9450 19932 10542
rect 20272 9586 20300 14758
rect 22112 11898 22140 19790
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 22756 14482 22784 17478
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 22744 14476 22796 14482
rect 22744 14418 22796 14424
rect 23664 14272 23716 14278
rect 23664 14214 23716 14220
rect 23676 12306 23704 14214
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 23664 12300 23716 12306
rect 23664 12242 23716 12248
rect 24676 12300 24728 12306
rect 24676 12242 24728 12248
rect 25412 12300 25464 12306
rect 25412 12242 25464 12248
rect 23296 12164 23348 12170
rect 23296 12106 23348 12112
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 21548 11824 21600 11830
rect 21548 11766 21600 11772
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20364 10130 20392 10406
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 20824 9994 20852 10542
rect 20916 10062 20944 11630
rect 20996 11280 21048 11286
rect 20996 11222 21048 11228
rect 20904 10056 20956 10062
rect 20904 9998 20956 10004
rect 20812 9988 20864 9994
rect 20812 9930 20864 9936
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 19892 9444 19944 9450
rect 19892 9386 19944 9392
rect 20168 9444 20220 9450
rect 20168 9386 20220 9392
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 19984 9104 20036 9110
rect 19984 9046 20036 9052
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 19444 8430 19472 8910
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 19444 7954 19472 8366
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19444 6390 19472 7346
rect 19904 7342 19932 7890
rect 19892 7336 19944 7342
rect 19892 7278 19944 7284
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 19432 6384 19484 6390
rect 19432 6326 19484 6332
rect 19904 6254 19932 7278
rect 19996 7206 20024 9046
rect 20076 9036 20128 9042
rect 20076 8978 20128 8984
rect 20088 8634 20116 8978
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 20180 8090 20208 9386
rect 20640 8838 20668 9522
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20260 8084 20312 8090
rect 20260 8026 20312 8032
rect 19984 7200 20036 7206
rect 19984 7142 20036 7148
rect 20168 6996 20220 7002
rect 20168 6938 20220 6944
rect 19892 6248 19944 6254
rect 19892 6190 19944 6196
rect 20180 6186 20208 6938
rect 20272 6934 20300 8026
rect 20536 7404 20588 7410
rect 20536 7346 20588 7352
rect 20444 7268 20496 7274
rect 20548 7256 20576 7346
rect 20496 7228 20576 7256
rect 20444 7210 20496 7216
rect 20260 6928 20312 6934
rect 20260 6870 20312 6876
rect 20732 6746 20760 9862
rect 20904 8832 20956 8838
rect 20904 8774 20956 8780
rect 20916 8362 20944 8774
rect 20904 8356 20956 8362
rect 20904 8298 20956 8304
rect 21008 7750 21036 11222
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 20996 7744 21048 7750
rect 20996 7686 21048 7692
rect 20640 6730 20760 6746
rect 20628 6724 20760 6730
rect 20680 6718 20760 6724
rect 20628 6666 20680 6672
rect 20168 6180 20220 6186
rect 20168 6122 20220 6128
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19352 5778 19380 6054
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 19340 5772 19392 5778
rect 19392 5732 19472 5760
rect 19340 5714 19392 5720
rect 19444 5234 19472 5732
rect 19432 5228 19484 5234
rect 19432 5170 19484 5176
rect 19444 4078 19472 5170
rect 20076 5092 20128 5098
rect 20076 5034 20128 5040
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 19892 4480 19944 4486
rect 19892 4422 19944 4428
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 19248 4004 19300 4010
rect 19248 3946 19300 3952
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19444 3194 19472 3470
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 19156 2984 19208 2990
rect 19156 2926 19208 2932
rect 16488 2916 16540 2922
rect 16488 2858 16540 2864
rect 16396 2848 16448 2854
rect 16396 2790 16448 2796
rect 18708 2582 18736 2926
rect 19904 2774 19932 4422
rect 19996 4282 20024 4422
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 20088 3194 20116 5034
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20628 4548 20680 4554
rect 20628 4490 20680 4496
rect 20444 4480 20496 4486
rect 20444 4422 20496 4428
rect 20456 4010 20484 4422
rect 20444 4004 20496 4010
rect 20444 3946 20496 3952
rect 20352 3392 20404 3398
rect 20352 3334 20404 3340
rect 20076 3188 20128 3194
rect 20076 3130 20128 3136
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19904 2746 20300 2774
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 15752 2576 15804 2582
rect 15752 2518 15804 2524
rect 18696 2576 18748 2582
rect 18696 2518 18748 2524
rect 20272 2446 20300 2746
rect 20364 2514 20392 3334
rect 20640 3058 20668 4490
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20732 2650 20760 4558
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 21100 2582 21128 9318
rect 21192 6662 21220 11018
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21284 8634 21312 10406
rect 21560 9110 21588 11766
rect 22112 9518 22140 11834
rect 22376 11688 22428 11694
rect 22376 11630 22428 11636
rect 22284 11008 22336 11014
rect 22284 10950 22336 10956
rect 22100 9512 22152 9518
rect 22100 9454 22152 9460
rect 21732 9376 21784 9382
rect 21732 9318 21784 9324
rect 21548 9104 21600 9110
rect 21548 9046 21600 9052
rect 21744 8974 21772 9318
rect 21732 8968 21784 8974
rect 21732 8910 21784 8916
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 21640 7200 21692 7206
rect 21640 7142 21692 7148
rect 21652 6934 21680 7142
rect 21640 6928 21692 6934
rect 21640 6870 21692 6876
rect 21180 6656 21232 6662
rect 21180 6598 21232 6604
rect 22204 6458 22232 8570
rect 22192 6452 22244 6458
rect 22192 6394 22244 6400
rect 21456 6248 21508 6254
rect 22192 6248 22244 6254
rect 21456 6190 21508 6196
rect 22190 6216 22192 6225
rect 22244 6216 22246 6225
rect 21468 6118 21496 6190
rect 21824 6180 21876 6186
rect 22296 6186 22324 10950
rect 22388 10606 22416 11630
rect 22468 11620 22520 11626
rect 22468 11562 22520 11568
rect 22376 10600 22428 10606
rect 22376 10542 22428 10548
rect 22388 9110 22416 10542
rect 22480 9654 22508 11562
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 23204 11144 23256 11150
rect 23204 11086 23256 11092
rect 22664 10810 22692 11086
rect 23216 11014 23244 11086
rect 23204 11008 23256 11014
rect 23204 10950 23256 10956
rect 22652 10804 22704 10810
rect 22652 10746 22704 10752
rect 22652 10532 22704 10538
rect 22652 10474 22704 10480
rect 22468 9648 22520 9654
rect 22468 9590 22520 9596
rect 22560 9512 22612 9518
rect 22560 9454 22612 9460
rect 22376 9104 22428 9110
rect 22376 9046 22428 9052
rect 22468 8968 22520 8974
rect 22572 8956 22600 9454
rect 22664 9382 22692 10474
rect 22744 10464 22796 10470
rect 22744 10406 22796 10412
rect 22756 9450 22784 10406
rect 23216 10062 23244 10950
rect 22928 10056 22980 10062
rect 22928 9998 22980 10004
rect 23204 10056 23256 10062
rect 23204 9998 23256 10004
rect 22744 9444 22796 9450
rect 22744 9386 22796 9392
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 22940 9178 22968 9998
rect 22928 9172 22980 9178
rect 22928 9114 22980 9120
rect 22520 8928 22600 8956
rect 22468 8910 22520 8916
rect 22572 8430 22600 8928
rect 22744 8968 22796 8974
rect 22744 8910 22796 8916
rect 22560 8424 22612 8430
rect 22560 8366 22612 8372
rect 22572 7886 22600 8366
rect 22560 7880 22612 7886
rect 22558 7848 22560 7857
rect 22612 7848 22614 7857
rect 22558 7783 22614 7792
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22388 6322 22416 7686
rect 22652 7268 22704 7274
rect 22652 7210 22704 7216
rect 22466 6896 22522 6905
rect 22466 6831 22522 6840
rect 22560 6860 22612 6866
rect 22480 6798 22508 6831
rect 22560 6802 22612 6808
rect 22468 6792 22520 6798
rect 22468 6734 22520 6740
rect 22376 6316 22428 6322
rect 22376 6258 22428 6264
rect 22572 6254 22600 6802
rect 22560 6248 22612 6254
rect 22560 6190 22612 6196
rect 22190 6151 22246 6160
rect 22284 6180 22336 6186
rect 21824 6122 21876 6128
rect 22284 6122 22336 6128
rect 21456 6112 21508 6118
rect 21456 6054 21508 6060
rect 21836 5930 21864 6122
rect 22100 6112 22152 6118
rect 22100 6054 22152 6060
rect 21560 5914 21864 5930
rect 21548 5908 21864 5914
rect 21600 5902 21864 5908
rect 21548 5850 21600 5856
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 21192 3194 21220 5170
rect 21456 3936 21508 3942
rect 21456 3878 21508 3884
rect 21180 3188 21232 3194
rect 21180 3130 21232 3136
rect 21468 2582 21496 3878
rect 21088 2576 21140 2582
rect 21088 2518 21140 2524
rect 21456 2576 21508 2582
rect 21456 2518 21508 2524
rect 20352 2508 20404 2514
rect 20352 2450 20404 2456
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 11060 2372 11112 2378
rect 11060 2314 11112 2320
rect 15568 2372 15620 2378
rect 15568 2314 15620 2320
rect 19984 2372 20036 2378
rect 19984 2314 20036 2320
rect 11072 800 11100 2314
rect 15580 800 15608 2314
rect 19996 800 20024 2314
rect 22112 2310 22140 6054
rect 22572 5794 22600 6190
rect 22480 5778 22600 5794
rect 22468 5772 22600 5778
rect 22520 5766 22600 5772
rect 22468 5714 22520 5720
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 22296 4146 22324 5646
rect 22572 5234 22600 5766
rect 22560 5228 22612 5234
rect 22560 5170 22612 5176
rect 22376 5024 22428 5030
rect 22376 4966 22428 4972
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 22388 3670 22416 4966
rect 22572 4690 22600 5170
rect 22560 4684 22612 4690
rect 22560 4626 22612 4632
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 22376 3664 22428 3670
rect 22376 3606 22428 3612
rect 22192 3596 22244 3602
rect 22192 3538 22244 3544
rect 22204 3058 22232 3538
rect 22480 3058 22508 3878
rect 22572 3602 22600 4626
rect 22664 3942 22692 7210
rect 22756 6730 22784 8910
rect 22928 8492 22980 8498
rect 22928 8434 22980 8440
rect 22940 8022 22968 8434
rect 22928 8016 22980 8022
rect 22928 7958 22980 7964
rect 22836 7880 22888 7886
rect 22836 7822 22888 7828
rect 22848 7546 22876 7822
rect 22836 7540 22888 7546
rect 22836 7482 22888 7488
rect 23308 6934 23336 12106
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 23400 11286 23428 12038
rect 23664 11688 23716 11694
rect 23664 11630 23716 11636
rect 23572 11552 23624 11558
rect 23572 11494 23624 11500
rect 23388 11280 23440 11286
rect 23388 11222 23440 11228
rect 23584 11218 23612 11494
rect 23676 11218 23704 11630
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 23572 11212 23624 11218
rect 23572 11154 23624 11160
rect 23664 11212 23716 11218
rect 23664 11154 23716 11160
rect 23584 10674 23612 11154
rect 23664 11076 23716 11082
rect 23664 11018 23716 11024
rect 23572 10668 23624 10674
rect 23572 10610 23624 10616
rect 23572 8356 23624 8362
rect 23572 8298 23624 8304
rect 23584 8090 23612 8298
rect 23480 8084 23532 8090
rect 23480 8026 23532 8032
rect 23572 8084 23624 8090
rect 23572 8026 23624 8032
rect 23492 7886 23520 8026
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 23676 7410 23704 11018
rect 23756 9988 23808 9994
rect 23756 9930 23808 9936
rect 23664 7404 23716 7410
rect 23664 7346 23716 7352
rect 23296 6928 23348 6934
rect 23296 6870 23348 6876
rect 22744 6724 22796 6730
rect 22744 6666 22796 6672
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 22848 5846 22876 6598
rect 23768 5846 23796 9930
rect 23848 9376 23900 9382
rect 23848 9318 23900 9324
rect 23860 6798 23888 9318
rect 24136 8242 24164 11494
rect 24400 11008 24452 11014
rect 24400 10950 24452 10956
rect 24412 10606 24440 10950
rect 24400 10600 24452 10606
rect 24400 10542 24452 10548
rect 24308 9580 24360 9586
rect 24308 9522 24360 9528
rect 24216 8832 24268 8838
rect 24216 8774 24268 8780
rect 24044 8214 24164 8242
rect 23848 6792 23900 6798
rect 23848 6734 23900 6740
rect 22836 5840 22888 5846
rect 22836 5782 22888 5788
rect 23756 5840 23808 5846
rect 23756 5782 23808 5788
rect 22836 5568 22888 5574
rect 22836 5510 22888 5516
rect 22848 4758 22876 5510
rect 24044 5166 24072 8214
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 24136 7002 24164 7482
rect 24228 7410 24256 8774
rect 24216 7404 24268 7410
rect 24216 7346 24268 7352
rect 24124 6996 24176 7002
rect 24124 6938 24176 6944
rect 24320 6458 24348 9522
rect 24412 6866 24440 10542
rect 24596 9110 24624 11494
rect 24688 10538 24716 12242
rect 25424 12102 25452 12242
rect 25412 12096 25464 12102
rect 25412 12038 25464 12044
rect 25424 11694 25452 12038
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 25228 11688 25280 11694
rect 25228 11630 25280 11636
rect 25412 11688 25464 11694
rect 25412 11630 25464 11636
rect 27988 11688 28040 11694
rect 27988 11630 28040 11636
rect 25240 11218 25268 11630
rect 25596 11620 25648 11626
rect 25596 11562 25648 11568
rect 25228 11212 25280 11218
rect 25228 11154 25280 11160
rect 24768 11144 24820 11150
rect 24768 11086 24820 11092
rect 24780 10606 24808 11086
rect 25608 10810 25636 11562
rect 26240 11144 26292 11150
rect 26240 11086 26292 11092
rect 25688 11076 25740 11082
rect 25688 11018 25740 11024
rect 25780 11076 25832 11082
rect 25780 11018 25832 11024
rect 25596 10804 25648 10810
rect 25596 10746 25648 10752
rect 24768 10600 24820 10606
rect 24768 10542 24820 10548
rect 24676 10532 24728 10538
rect 24676 10474 24728 10480
rect 24688 10130 24716 10474
rect 24780 10130 24808 10542
rect 24676 10124 24728 10130
rect 24676 10066 24728 10072
rect 24768 10124 24820 10130
rect 24768 10066 24820 10072
rect 25228 10056 25280 10062
rect 25228 9998 25280 10004
rect 24860 9920 24912 9926
rect 24860 9862 24912 9868
rect 24676 9172 24728 9178
rect 24676 9114 24728 9120
rect 24584 9104 24636 9110
rect 24584 9046 24636 9052
rect 24490 7848 24546 7857
rect 24490 7783 24546 7792
rect 24504 7410 24532 7783
rect 24492 7404 24544 7410
rect 24492 7346 24544 7352
rect 24400 6860 24452 6866
rect 24400 6802 24452 6808
rect 24308 6452 24360 6458
rect 24308 6394 24360 6400
rect 24124 5908 24176 5914
rect 24124 5850 24176 5856
rect 24136 5574 24164 5850
rect 24412 5778 24440 6802
rect 24400 5772 24452 5778
rect 24400 5714 24452 5720
rect 24124 5568 24176 5574
rect 24124 5510 24176 5516
rect 24032 5160 24084 5166
rect 24032 5102 24084 5108
rect 22836 4752 22888 4758
rect 22836 4694 22888 4700
rect 22928 4276 22980 4282
rect 22928 4218 22980 4224
rect 22836 4004 22888 4010
rect 22836 3946 22888 3952
rect 22652 3936 22704 3942
rect 22652 3878 22704 3884
rect 22560 3596 22612 3602
rect 22560 3538 22612 3544
rect 22848 3398 22876 3946
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22192 3052 22244 3058
rect 22192 2994 22244 3000
rect 22468 3052 22520 3058
rect 22468 2994 22520 3000
rect 22204 2774 22232 2994
rect 22204 2746 22324 2774
rect 22296 2514 22324 2746
rect 22940 2650 22968 4218
rect 23112 4208 23164 4214
rect 23112 4150 23164 4156
rect 23124 2650 23152 4150
rect 23664 4004 23716 4010
rect 23664 3946 23716 3952
rect 24216 4004 24268 4010
rect 24216 3946 24268 3952
rect 23676 3641 23704 3946
rect 24228 3738 24256 3946
rect 24216 3732 24268 3738
rect 24216 3674 24268 3680
rect 24584 3732 24636 3738
rect 24584 3674 24636 3680
rect 23662 3632 23718 3641
rect 23662 3567 23718 3576
rect 24596 2922 24624 3674
rect 24688 2990 24716 9114
rect 24872 8634 24900 9862
rect 25240 9586 25268 9998
rect 25228 9580 25280 9586
rect 25228 9522 25280 9528
rect 25134 9480 25190 9489
rect 24952 9444 25004 9450
rect 25134 9415 25190 9424
rect 24952 9386 25004 9392
rect 24964 9178 24992 9386
rect 24952 9172 25004 9178
rect 24952 9114 25004 9120
rect 25148 9042 25176 9415
rect 25136 9036 25188 9042
rect 25136 8978 25188 8984
rect 25042 8664 25098 8673
rect 24860 8628 24912 8634
rect 25042 8599 25098 8608
rect 24860 8570 24912 8576
rect 25056 8362 25084 8599
rect 25044 8356 25096 8362
rect 25044 8298 25096 8304
rect 25148 7886 25176 8978
rect 25240 8430 25268 9522
rect 25504 9376 25556 9382
rect 25504 9318 25556 9324
rect 25596 9376 25648 9382
rect 25596 9318 25648 9324
rect 25516 9110 25544 9318
rect 25504 9104 25556 9110
rect 25504 9046 25556 9052
rect 25608 8566 25636 9318
rect 25596 8560 25648 8566
rect 25596 8502 25648 8508
rect 25228 8424 25280 8430
rect 25228 8366 25280 8372
rect 25320 8288 25372 8294
rect 25320 8230 25372 8236
rect 25332 8106 25360 8230
rect 25332 8078 25636 8106
rect 25608 7886 25636 8078
rect 25136 7880 25188 7886
rect 25136 7822 25188 7828
rect 25504 7880 25556 7886
rect 25504 7822 25556 7828
rect 25596 7880 25648 7886
rect 25596 7822 25648 7828
rect 24952 7744 25004 7750
rect 24952 7686 25004 7692
rect 24964 7546 24992 7686
rect 24952 7540 25004 7546
rect 24952 7482 25004 7488
rect 25320 7540 25372 7546
rect 25320 7482 25372 7488
rect 25332 6934 25360 7482
rect 25412 7404 25464 7410
rect 25412 7346 25464 7352
rect 25320 6928 25372 6934
rect 25320 6870 25372 6876
rect 24952 6792 25004 6798
rect 24952 6734 25004 6740
rect 24860 6452 24912 6458
rect 24860 6394 24912 6400
rect 24872 6254 24900 6394
rect 24860 6248 24912 6254
rect 24860 6190 24912 6196
rect 24768 6112 24820 6118
rect 24768 6054 24820 6060
rect 24780 5234 24808 6054
rect 24860 5840 24912 5846
rect 24860 5782 24912 5788
rect 24872 5370 24900 5782
rect 24860 5364 24912 5370
rect 24860 5306 24912 5312
rect 24964 5302 24992 6734
rect 25226 6080 25282 6089
rect 25226 6015 25282 6024
rect 25240 5778 25268 6015
rect 25424 5914 25452 7346
rect 25516 6905 25544 7822
rect 25700 6934 25728 11018
rect 25792 10266 25820 11018
rect 26148 11008 26200 11014
rect 26148 10950 26200 10956
rect 25964 10464 26016 10470
rect 25964 10406 26016 10412
rect 25780 10260 25832 10266
rect 25780 10202 25832 10208
rect 25792 10062 25820 10202
rect 25780 10056 25832 10062
rect 25780 9998 25832 10004
rect 25780 9444 25832 9450
rect 25780 9386 25832 9392
rect 25792 8634 25820 9386
rect 25780 8628 25832 8634
rect 25780 8570 25832 8576
rect 25780 8288 25832 8294
rect 25780 8230 25832 8236
rect 25792 8022 25820 8230
rect 25780 8016 25832 8022
rect 25780 7958 25832 7964
rect 25976 7274 26004 10406
rect 26160 10130 26188 10950
rect 26252 10606 26280 11086
rect 27068 10668 27120 10674
rect 27068 10610 27120 10616
rect 26240 10600 26292 10606
rect 26240 10542 26292 10548
rect 26252 10130 26280 10542
rect 26148 10124 26200 10130
rect 26148 10066 26200 10072
rect 26240 10124 26292 10130
rect 26240 10066 26292 10072
rect 26160 9081 26188 10066
rect 26516 9512 26568 9518
rect 26514 9480 26516 9489
rect 26568 9480 26570 9489
rect 26240 9444 26292 9450
rect 26570 9438 26740 9466
rect 26514 9415 26570 9424
rect 26240 9386 26292 9392
rect 26146 9072 26202 9081
rect 26146 9007 26202 9016
rect 26252 8090 26280 9386
rect 26516 9104 26568 9110
rect 26516 9046 26568 9052
rect 26528 8634 26556 9046
rect 26608 8832 26660 8838
rect 26608 8774 26660 8780
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 26240 8084 26292 8090
rect 26240 8026 26292 8032
rect 26620 7750 26648 8774
rect 26712 8344 26740 9438
rect 26792 8356 26844 8362
rect 26712 8316 26792 8344
rect 26608 7744 26660 7750
rect 26608 7686 26660 7692
rect 26712 7410 26740 8316
rect 26792 8298 26844 8304
rect 26792 7744 26844 7750
rect 26792 7686 26844 7692
rect 26700 7404 26752 7410
rect 26700 7346 26752 7352
rect 25964 7268 26016 7274
rect 25964 7210 26016 7216
rect 26712 6934 26740 7346
rect 25688 6928 25740 6934
rect 25502 6896 25558 6905
rect 25688 6870 25740 6876
rect 26700 6928 26752 6934
rect 26700 6870 26752 6876
rect 25502 6831 25558 6840
rect 26148 6656 26200 6662
rect 26148 6598 26200 6604
rect 26160 6186 26188 6598
rect 26516 6248 26568 6254
rect 26422 6216 26478 6225
rect 26148 6180 26200 6186
rect 26516 6190 26568 6196
rect 26422 6151 26478 6160
rect 26148 6122 26200 6128
rect 25412 5908 25464 5914
rect 25412 5850 25464 5856
rect 25228 5772 25280 5778
rect 25228 5714 25280 5720
rect 24952 5296 25004 5302
rect 24952 5238 25004 5244
rect 24768 5228 24820 5234
rect 24768 5170 24820 5176
rect 24860 4140 24912 4146
rect 24860 4082 24912 4088
rect 24872 3602 24900 4082
rect 25240 4010 25268 5714
rect 25872 5228 25924 5234
rect 25872 5170 25924 5176
rect 25884 4758 25912 5170
rect 26332 5092 26384 5098
rect 26332 5034 26384 5040
rect 25872 4752 25924 4758
rect 25872 4694 25924 4700
rect 26240 4752 26292 4758
rect 26240 4694 26292 4700
rect 25228 4004 25280 4010
rect 25228 3946 25280 3952
rect 25240 3602 25268 3946
rect 24860 3596 24912 3602
rect 24860 3538 24912 3544
rect 25228 3596 25280 3602
rect 25228 3538 25280 3544
rect 24676 2984 24728 2990
rect 24676 2926 24728 2932
rect 24584 2916 24636 2922
rect 24584 2858 24636 2864
rect 25044 2848 25096 2854
rect 25044 2790 25096 2796
rect 22928 2644 22980 2650
rect 22928 2586 22980 2592
rect 23112 2644 23164 2650
rect 23112 2586 23164 2592
rect 25056 2582 25084 2790
rect 25044 2576 25096 2582
rect 25044 2518 25096 2524
rect 25240 2514 25268 3538
rect 26252 3126 26280 4694
rect 26344 3194 26372 5034
rect 26332 3188 26384 3194
rect 26332 3130 26384 3136
rect 26240 3120 26292 3126
rect 26240 3062 26292 3068
rect 25780 2984 25832 2990
rect 25780 2926 25832 2932
rect 25792 2650 25820 2926
rect 26436 2774 26464 6151
rect 26528 6089 26556 6190
rect 26514 6080 26570 6089
rect 26514 6015 26570 6024
rect 26712 5234 26740 6870
rect 26804 6458 26832 7686
rect 26792 6452 26844 6458
rect 26792 6394 26844 6400
rect 26976 6180 27028 6186
rect 26976 6122 27028 6128
rect 26988 5914 27016 6122
rect 26976 5908 27028 5914
rect 26976 5850 27028 5856
rect 26700 5228 26752 5234
rect 26752 5188 26832 5216
rect 26700 5170 26752 5176
rect 26804 4622 26832 5188
rect 26700 4616 26752 4622
rect 26700 4558 26752 4564
rect 26792 4616 26844 4622
rect 26792 4558 26844 4564
rect 26712 4486 26740 4558
rect 26608 4480 26660 4486
rect 26608 4422 26660 4428
rect 26700 4480 26752 4486
rect 26700 4422 26752 4428
rect 26620 3194 26648 4422
rect 26700 3936 26752 3942
rect 26700 3878 26752 3884
rect 26608 3188 26660 3194
rect 26608 3130 26660 3136
rect 26712 2990 26740 3878
rect 27080 3738 27108 10610
rect 27160 10124 27212 10130
rect 27160 10066 27212 10072
rect 27344 10124 27396 10130
rect 27344 10066 27396 10072
rect 27172 10010 27200 10066
rect 27172 9982 27292 10010
rect 27160 9920 27212 9926
rect 27160 9862 27212 9868
rect 27172 7206 27200 9862
rect 27160 7200 27212 7206
rect 27160 7142 27212 7148
rect 27264 6730 27292 9982
rect 27356 9586 27384 10066
rect 27804 9648 27856 9654
rect 27804 9590 27856 9596
rect 27344 9580 27396 9586
rect 27344 9522 27396 9528
rect 27618 9072 27674 9081
rect 27618 9007 27620 9016
rect 27672 9007 27674 9016
rect 27620 8978 27672 8984
rect 27712 8900 27764 8906
rect 27712 8842 27764 8848
rect 27344 8424 27396 8430
rect 27344 8366 27396 8372
rect 27356 7954 27384 8366
rect 27344 7948 27396 7954
rect 27344 7890 27396 7896
rect 27252 6724 27304 6730
rect 27252 6666 27304 6672
rect 27356 6633 27384 7890
rect 27724 7410 27752 8842
rect 27712 7404 27764 7410
rect 27712 7346 27764 7352
rect 27816 6934 27844 9590
rect 28000 9518 28028 11630
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 30012 10804 30064 10810
rect 30012 10746 30064 10752
rect 27988 9512 28040 9518
rect 27988 9454 28040 9460
rect 28908 9444 28960 9450
rect 28908 9386 28960 9392
rect 28448 9376 28500 9382
rect 28448 9318 28500 9324
rect 28460 8673 28488 9318
rect 28920 9042 28948 9386
rect 28908 9036 28960 9042
rect 28908 8978 28960 8984
rect 28446 8664 28502 8673
rect 28446 8599 28502 8608
rect 28920 7886 28948 8978
rect 29184 8424 29236 8430
rect 29184 8366 29236 8372
rect 28908 7880 28960 7886
rect 28908 7822 28960 7828
rect 29196 7546 29224 8366
rect 29552 8288 29604 8294
rect 29552 8230 29604 8236
rect 29564 8022 29592 8230
rect 29552 8016 29604 8022
rect 29552 7958 29604 7964
rect 29276 7948 29328 7954
rect 29276 7890 29328 7896
rect 28632 7540 28684 7546
rect 28632 7482 28684 7488
rect 29184 7540 29236 7546
rect 29184 7482 29236 7488
rect 28172 7404 28224 7410
rect 28172 7346 28224 7352
rect 28184 7274 28212 7346
rect 28172 7268 28224 7274
rect 28172 7210 28224 7216
rect 27804 6928 27856 6934
rect 27804 6870 27856 6876
rect 27436 6860 27488 6866
rect 27436 6802 27488 6808
rect 27342 6624 27398 6633
rect 27342 6559 27398 6568
rect 27252 6452 27304 6458
rect 27252 6394 27304 6400
rect 27068 3732 27120 3738
rect 27068 3674 27120 3680
rect 27264 3602 27292 6394
rect 27356 3602 27384 6559
rect 27448 6254 27476 6802
rect 27436 6248 27488 6254
rect 27436 6190 27488 6196
rect 28172 6112 28224 6118
rect 28172 6054 28224 6060
rect 28184 5710 28212 6054
rect 28448 5840 28500 5846
rect 28448 5782 28500 5788
rect 28172 5704 28224 5710
rect 28172 5646 28224 5652
rect 28356 5704 28408 5710
rect 28356 5646 28408 5652
rect 27436 5568 27488 5574
rect 28172 5568 28224 5574
rect 27436 5510 27488 5516
rect 28170 5536 28172 5545
rect 28264 5568 28316 5574
rect 28224 5536 28226 5545
rect 27448 4282 27476 5510
rect 28264 5510 28316 5516
rect 28170 5471 28226 5480
rect 28276 5302 28304 5510
rect 28264 5296 28316 5302
rect 28264 5238 28316 5244
rect 27988 5092 28040 5098
rect 27988 5034 28040 5040
rect 27896 5024 27948 5030
rect 27896 4966 27948 4972
rect 27804 4684 27856 4690
rect 27804 4626 27856 4632
rect 27816 4282 27844 4626
rect 27436 4276 27488 4282
rect 27436 4218 27488 4224
rect 27804 4276 27856 4282
rect 27804 4218 27856 4224
rect 27908 4146 27936 4966
rect 27620 4140 27672 4146
rect 27620 4082 27672 4088
rect 27896 4140 27948 4146
rect 27896 4082 27948 4088
rect 27632 3738 27660 4082
rect 27896 4004 27948 4010
rect 27896 3946 27948 3952
rect 27620 3732 27672 3738
rect 27620 3674 27672 3680
rect 27252 3596 27304 3602
rect 27252 3538 27304 3544
rect 27344 3596 27396 3602
rect 27344 3538 27396 3544
rect 27908 3534 27936 3946
rect 26792 3528 26844 3534
rect 26792 3470 26844 3476
rect 27896 3528 27948 3534
rect 27896 3470 27948 3476
rect 26700 2984 26752 2990
rect 26700 2926 26752 2932
rect 26436 2746 26648 2774
rect 26620 2650 26648 2746
rect 25780 2644 25832 2650
rect 25780 2586 25832 2592
rect 26608 2644 26660 2650
rect 26608 2586 26660 2592
rect 26804 2514 26832 3470
rect 28000 3466 28028 5034
rect 28264 4616 28316 4622
rect 28264 4558 28316 4564
rect 28172 4072 28224 4078
rect 28172 4014 28224 4020
rect 28184 3602 28212 4014
rect 28276 4010 28304 4558
rect 28368 4486 28396 5646
rect 28356 4480 28408 4486
rect 28356 4422 28408 4428
rect 28264 4004 28316 4010
rect 28264 3946 28316 3952
rect 28172 3596 28224 3602
rect 28172 3538 28224 3544
rect 28184 3482 28212 3538
rect 27988 3460 28040 3466
rect 27988 3402 28040 3408
rect 28092 3454 28212 3482
rect 26884 3188 26936 3194
rect 26884 3130 26936 3136
rect 26976 3188 27028 3194
rect 26976 3130 27028 3136
rect 26896 2650 26924 3130
rect 26884 2644 26936 2650
rect 26884 2586 26936 2592
rect 26988 2582 27016 3130
rect 27068 3120 27120 3126
rect 27068 3062 27120 3068
rect 26976 2576 27028 2582
rect 26976 2518 27028 2524
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 25228 2508 25280 2514
rect 25228 2450 25280 2456
rect 26792 2508 26844 2514
rect 26792 2450 26844 2456
rect 27080 2378 27108 3062
rect 28092 2774 28120 3454
rect 28276 2922 28304 3946
rect 28354 3632 28410 3641
rect 28354 3567 28410 3576
rect 28368 3534 28396 3567
rect 28356 3528 28408 3534
rect 28356 3470 28408 3476
rect 28356 2984 28408 2990
rect 28356 2926 28408 2932
rect 28264 2916 28316 2922
rect 28264 2858 28316 2864
rect 28092 2746 28212 2774
rect 28184 2446 28212 2746
rect 28276 2650 28304 2858
rect 28368 2666 28396 2926
rect 28460 2854 28488 5782
rect 28644 3942 28672 7482
rect 29288 7410 29316 7890
rect 29276 7404 29328 7410
rect 29276 7346 29328 7352
rect 29552 7404 29604 7410
rect 29552 7346 29604 7352
rect 28724 7200 28776 7206
rect 28724 7142 28776 7148
rect 28736 4758 28764 7142
rect 28816 6656 28868 6662
rect 28814 6624 28816 6633
rect 29368 6656 29420 6662
rect 28868 6624 28870 6633
rect 29368 6598 29420 6604
rect 28814 6559 28870 6568
rect 29380 6254 29408 6598
rect 29368 6248 29420 6254
rect 29368 6190 29420 6196
rect 28814 6080 28870 6089
rect 28814 6015 28870 6024
rect 28828 5846 28856 6015
rect 28816 5840 28868 5846
rect 28816 5782 28868 5788
rect 29276 5772 29328 5778
rect 29276 5714 29328 5720
rect 29288 5658 29316 5714
rect 29196 5630 29316 5658
rect 29368 5636 29420 5642
rect 28908 5024 28960 5030
rect 28908 4966 28960 4972
rect 28724 4752 28776 4758
rect 28724 4694 28776 4700
rect 28632 3936 28684 3942
rect 28632 3878 28684 3884
rect 28920 3602 28948 4966
rect 29196 4690 29224 5630
rect 29368 5578 29420 5584
rect 29276 5092 29328 5098
rect 29276 5034 29328 5040
rect 29288 4826 29316 5034
rect 29276 4820 29328 4826
rect 29276 4762 29328 4768
rect 29184 4684 29236 4690
rect 29184 4626 29236 4632
rect 29000 3936 29052 3942
rect 29000 3878 29052 3884
rect 29012 3670 29040 3878
rect 29000 3664 29052 3670
rect 29000 3606 29052 3612
rect 28540 3596 28592 3602
rect 28540 3538 28592 3544
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 28448 2848 28500 2854
rect 28448 2790 28500 2796
rect 28552 2666 28580 3538
rect 29196 3194 29224 4626
rect 29380 4078 29408 5578
rect 29564 5166 29592 7346
rect 30024 7342 30052 10746
rect 31300 9920 31352 9926
rect 31300 9862 31352 9868
rect 30380 9512 30432 9518
rect 30380 9454 30432 9460
rect 30196 8968 30248 8974
rect 30196 8910 30248 8916
rect 30208 7478 30236 8910
rect 30392 8430 30420 9454
rect 30472 9104 30524 9110
rect 30472 9046 30524 9052
rect 30380 8424 30432 8430
rect 30380 8366 30432 8372
rect 30288 8084 30340 8090
rect 30288 8026 30340 8032
rect 30196 7472 30248 7478
rect 30196 7414 30248 7420
rect 30012 7336 30064 7342
rect 30012 7278 30064 7284
rect 29828 7268 29880 7274
rect 29828 7210 29880 7216
rect 29840 6458 29868 7210
rect 30024 6934 30052 7278
rect 30012 6928 30064 6934
rect 30012 6870 30064 6876
rect 29828 6452 29880 6458
rect 29828 6394 29880 6400
rect 30024 5710 30052 6870
rect 30208 6338 30236 7414
rect 30300 6458 30328 8026
rect 30380 7200 30432 7206
rect 30380 7142 30432 7148
rect 30288 6452 30340 6458
rect 30288 6394 30340 6400
rect 30208 6310 30328 6338
rect 30300 6254 30328 6310
rect 30288 6248 30340 6254
rect 30288 6190 30340 6196
rect 30012 5704 30064 5710
rect 30012 5646 30064 5652
rect 30024 5166 30052 5646
rect 30300 5642 30328 6190
rect 30392 5914 30420 7142
rect 30484 6866 30512 9046
rect 31312 7954 31340 9862
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 31484 8424 31536 8430
rect 31484 8366 31536 8372
rect 31300 7948 31352 7954
rect 31300 7890 31352 7896
rect 30840 7336 30892 7342
rect 30840 7278 30892 7284
rect 30472 6860 30524 6866
rect 30472 6802 30524 6808
rect 30852 6662 30880 7278
rect 31312 6934 31340 7890
rect 31496 7342 31524 8366
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 31484 7336 31536 7342
rect 31484 7278 31536 7284
rect 31300 6928 31352 6934
rect 31300 6870 31352 6876
rect 30840 6656 30892 6662
rect 30840 6598 30892 6604
rect 31668 6656 31720 6662
rect 31668 6598 31720 6604
rect 32404 6656 32456 6662
rect 32404 6598 32456 6604
rect 30472 6384 30524 6390
rect 30472 6326 30524 6332
rect 30380 5908 30432 5914
rect 30380 5850 30432 5856
rect 30288 5636 30340 5642
rect 30288 5578 30340 5584
rect 30484 5574 30512 6326
rect 31680 6186 31708 6598
rect 31668 6180 31720 6186
rect 31668 6122 31720 6128
rect 31680 5846 31708 6122
rect 31944 6112 31996 6118
rect 31944 6054 31996 6060
rect 31392 5840 31444 5846
rect 31392 5782 31444 5788
rect 31668 5840 31720 5846
rect 31668 5782 31720 5788
rect 31300 5772 31352 5778
rect 31300 5714 31352 5720
rect 31312 5574 31340 5714
rect 30472 5568 30524 5574
rect 30378 5536 30434 5545
rect 30472 5510 30524 5516
rect 31300 5568 31352 5574
rect 31300 5510 31352 5516
rect 30378 5471 30434 5480
rect 30392 5302 30420 5471
rect 30380 5296 30432 5302
rect 30380 5238 30432 5244
rect 31312 5166 31340 5510
rect 29552 5160 29604 5166
rect 29552 5102 29604 5108
rect 30012 5160 30064 5166
rect 30012 5102 30064 5108
rect 30656 5160 30708 5166
rect 30656 5102 30708 5108
rect 31300 5160 31352 5166
rect 31300 5102 31352 5108
rect 30668 4690 30696 5102
rect 30656 4684 30708 4690
rect 30656 4626 30708 4632
rect 30472 4480 30524 4486
rect 30472 4422 30524 4428
rect 30484 4214 30512 4422
rect 30472 4208 30524 4214
rect 30472 4150 30524 4156
rect 30668 4146 30696 4626
rect 30656 4140 30708 4146
rect 30656 4082 30708 4088
rect 29368 4072 29420 4078
rect 29368 4014 29420 4020
rect 29644 3936 29696 3942
rect 29644 3878 29696 3884
rect 29552 3596 29604 3602
rect 29552 3538 29604 3544
rect 29184 3188 29236 3194
rect 29184 3130 29236 3136
rect 29564 2990 29592 3538
rect 29656 3058 29684 3878
rect 31404 3602 31432 5782
rect 31760 5568 31812 5574
rect 31760 5510 31812 5516
rect 31392 3596 31444 3602
rect 31392 3538 31444 3544
rect 31772 3466 31800 5510
rect 31956 5234 31984 6054
rect 32416 5710 32444 6598
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 32404 5704 32456 5710
rect 32404 5646 32456 5652
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 31944 5228 31996 5234
rect 31944 5170 31996 5176
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 31760 3460 31812 3466
rect 31760 3402 31812 3408
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 29644 3052 29696 3058
rect 29644 2994 29696 3000
rect 29552 2984 29604 2990
rect 29552 2926 29604 2932
rect 28724 2916 28776 2922
rect 28724 2858 28776 2864
rect 28264 2644 28316 2650
rect 28264 2586 28316 2592
rect 28368 2638 28580 2666
rect 28368 2514 28396 2638
rect 28356 2508 28408 2514
rect 28356 2450 28408 2456
rect 28172 2440 28224 2446
rect 28172 2382 28224 2388
rect 27068 2372 27120 2378
rect 27068 2314 27120 2320
rect 22100 2304 22152 2310
rect 22100 2246 22152 2252
rect 28736 1018 28764 2858
rect 28908 2372 28960 2378
rect 28908 2314 28960 2320
rect 33324 2372 33376 2378
rect 33324 2314 33376 2320
rect 37740 2372 37792 2378
rect 37740 2314 37792 2320
rect 24400 1012 24452 1018
rect 24400 954 24452 960
rect 28724 1012 28776 1018
rect 28724 954 28776 960
rect 24412 800 24440 954
rect 28920 800 28948 2314
rect 33336 800 33364 2314
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 37752 800 37780 2314
rect 2226 0 2282 800
rect 6642 0 6698 800
rect 11058 0 11114 800
rect 15566 0 15622 800
rect 19982 0 20038 800
rect 24398 0 24454 800
rect 28906 0 28962 800
rect 33322 0 33378 800
rect 37738 0 37794 800
<< via2 >>
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 22190 6196 22192 6216
rect 22192 6196 22244 6216
rect 22244 6196 22246 6216
rect 22190 6160 22246 6196
rect 22558 7828 22560 7848
rect 22560 7828 22612 7848
rect 22612 7828 22614 7848
rect 22558 7792 22614 7828
rect 22466 6840 22522 6896
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 24490 7792 24546 7848
rect 23662 3576 23718 3632
rect 25134 9424 25190 9480
rect 25042 8608 25098 8664
rect 25226 6024 25282 6080
rect 26514 9460 26516 9480
rect 26516 9460 26568 9480
rect 26568 9460 26570 9480
rect 26514 9424 26570 9460
rect 26146 9016 26202 9072
rect 25502 6840 25558 6896
rect 26422 6160 26478 6216
rect 26514 6024 26570 6080
rect 27618 9036 27674 9072
rect 27618 9016 27620 9036
rect 27620 9016 27672 9036
rect 27672 9016 27674 9036
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 28446 8608 28502 8664
rect 27342 6568 27398 6624
rect 28170 5516 28172 5536
rect 28172 5516 28224 5536
rect 28224 5516 28226 5536
rect 28170 5480 28226 5516
rect 28354 3576 28410 3632
rect 28814 6604 28816 6624
rect 28816 6604 28868 6624
rect 28868 6604 28870 6624
rect 28814 6568 28870 6604
rect 28814 6024 28870 6080
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 30378 5480 30434 5536
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
<< metal3 >>
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 28255 35248 28256
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 27167 35248 27168
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 16287 35248 16288
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 13023 35248 13024
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 10847 35248 10848
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 25129 9482 25195 9485
rect 26509 9482 26575 9485
rect 25129 9480 26575 9482
rect 25129 9424 25134 9480
rect 25190 9424 26514 9480
rect 26570 9424 26575 9480
rect 25129 9422 26575 9424
rect 25129 9419 25195 9422
rect 26509 9419 26575 9422
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 26141 9074 26207 9077
rect 27613 9074 27679 9077
rect 26141 9072 27679 9074
rect 26141 9016 26146 9072
rect 26202 9016 27618 9072
rect 27674 9016 27679 9072
rect 26141 9014 27679 9016
rect 26141 9011 26207 9014
rect 27613 9011 27679 9014
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 25037 8666 25103 8669
rect 28441 8666 28507 8669
rect 25037 8664 28507 8666
rect 25037 8608 25042 8664
rect 25098 8608 28446 8664
rect 28502 8608 28507 8664
rect 25037 8606 28507 8608
rect 25037 8603 25103 8606
rect 28441 8603 28507 8606
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 22553 7850 22619 7853
rect 24485 7850 24551 7853
rect 22553 7848 24551 7850
rect 22553 7792 22558 7848
rect 22614 7792 24490 7848
rect 24546 7792 24551 7848
rect 22553 7790 24551 7792
rect 22553 7787 22619 7790
rect 24485 7787 24551 7790
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 22461 6898 22527 6901
rect 25497 6898 25563 6901
rect 22461 6896 25563 6898
rect 22461 6840 22466 6896
rect 22522 6840 25502 6896
rect 25558 6840 25563 6896
rect 22461 6838 25563 6840
rect 22461 6835 22527 6838
rect 25497 6835 25563 6838
rect 27337 6626 27403 6629
rect 28809 6626 28875 6629
rect 27337 6624 28875 6626
rect 27337 6568 27342 6624
rect 27398 6568 28814 6624
rect 28870 6568 28875 6624
rect 27337 6566 28875 6568
rect 27337 6563 27403 6566
rect 28809 6563 28875 6566
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 6495 35248 6496
rect 22185 6218 22251 6221
rect 26417 6218 26483 6221
rect 22185 6216 26483 6218
rect 22185 6160 22190 6216
rect 22246 6160 26422 6216
rect 26478 6160 26483 6216
rect 22185 6158 26483 6160
rect 22185 6155 22251 6158
rect 26417 6155 26483 6158
rect 25221 6082 25287 6085
rect 26509 6082 26575 6085
rect 28809 6082 28875 6085
rect 25221 6080 28875 6082
rect 25221 6024 25226 6080
rect 25282 6024 26514 6080
rect 26570 6024 28814 6080
rect 28870 6024 28875 6080
rect 25221 6022 28875 6024
rect 25221 6019 25287 6022
rect 26509 6019 26575 6022
rect 28809 6019 28875 6022
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 28165 5538 28231 5541
rect 30373 5538 30439 5541
rect 28165 5536 30439 5538
rect 28165 5480 28170 5536
rect 28226 5480 30378 5536
rect 30434 5480 30439 5536
rect 28165 5478 30439 5480
rect 28165 5475 28231 5478
rect 30373 5475 30439 5478
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 23657 3634 23723 3637
rect 28349 3634 28415 3637
rect 23657 3632 28415 3634
rect 23657 3576 23662 3632
rect 23718 3576 28354 3632
rect 28410 3576 28415 3632
rect 23657 3574 28415 3576
rect 23657 3571 23723 3574
rect 28349 3571 28415 3574
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
<< via3 >>
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
<< metal4 >>
rect 4208 37024 4528 37584
rect 19568 37568 19888 37584
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4868 2176 5188 37536
rect 5528 2176 5848 37536
rect 6188 2176 6508 37536
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 4208 2128 4528 2144
rect 19568 2128 19888 2688
rect 20228 2176 20548 37536
rect 20888 2176 21208 37536
rect 21548 2176 21868 37536
rect 34928 37024 35248 37584
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 35588 2176 35908 37536
rect 36248 2176 36568 37536
rect 36908 2176 37228 37536
rect 34928 2128 35248 2144
use sky130_fd_sc_hd__conb_1  _181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 2944 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1623529830
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform -1 0 2576 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 1380 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 2116 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 2576 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1623529830
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 3220 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_30
timestamp 1623529830
transform 1 0 3864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_42
timestamp 1623529830
transform 1 0 4968 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1623529830
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1623529830
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1623529830
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1623529830
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54
timestamp 1623529830
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_59
timestamp 1623529830
transform 1 0 6532 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_51
timestamp 1623529830
transform 1 0 5796 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_58
timestamp 1623529830
transform 1 0 6440 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1623529830
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_71
timestamp 1623529830
transform 1 0 7636 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1623529830
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_70
timestamp 1623529830
transform 1 0 7544 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_82
timestamp 1623529830
transform 1 0 8648 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _180_
timestamp 1623529830
transform -1 0 11224 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output8
timestamp 1623529830
transform -1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_88
timestamp 1623529830
transform 1 0 9200 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100
timestamp 1623529830
transform 1 0 10304 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_94
timestamp 1623529830
transform 1 0 9752 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_106
timestamp 1623529830
transform 1 0 10856 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1623529830
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1623529830
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1623529830
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_117
timestamp 1623529830
transform 1 0 11868 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_129
timestamp 1623529830
transform 1 0 12972 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_110
timestamp 1623529830
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_115
timestamp 1623529830
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_127
timestamp 1623529830
transform 1 0 12788 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1623529830
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1623529830
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_146
timestamp 1623529830
transform 1 0 14536 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_139
timestamp 1623529830
transform 1 0 13892 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_151
timestamp 1623529830
transform 1 0 14996 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _184_
timestamp 1623529830
transform 1 0 16468 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1623529830
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1623529830
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output3
timestamp 1623529830
transform -1 0 15916 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_154
timestamp 1623529830
transform 1 0 15272 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1623529830
transform 1 0 15916 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_170
timestamp 1623529830
transform 1 0 16744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_163
timestamp 1623529830
transform 1 0 16100 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_172
timestamp 1623529830
transform 1 0 16928 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform -1 0 18400 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform -1 0 19504 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _172_
timestamp 1623529830
transform -1 0 19412 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output7
timestamp 1623529830
transform 1 0 17940 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_175
timestamp 1623529830
transform 1 0 17204 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1623529830
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_180
timestamp 1623529830
transform 1 0 17664 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1623529830
transform 1 0 18400 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _228_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform -1 0 21712 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _230_
timestamp 1623529830
transform -1 0 22080 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1623529830
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_199
timestamp 1623529830
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_204
timestamp 1623529830
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_200
timestamp 1623529830
transform 1 0 19504 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _207_
timestamp 1623529830
transform 1 0 22540 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _209_
timestamp 1623529830
transform -1 0 24748 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1623529830
transform 1 0 22448 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1623529830
transform 1 0 22080 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_228
timestamp 1623529830
transform 1 0 22080 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_233
timestamp 1623529830
transform 1 0 22540 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_224
timestamp 1623529830
transform 1 0 21712 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_229
timestamp 1623529830
transform 1 0 22172 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 24748 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1623529830
transform 1 0 25116 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_257
timestamp 1623529830
transform 1 0 24748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1623529830
transform 1 0 25208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_253
timestamp 1623529830
transform 1 0 24380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_260
timestamp 1623529830
transform 1 0 25024 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_267
timestamp 1623529830
transform 1 0 25668 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_269
timestamp 1623529830
transform 1 0 25852 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1623529830
transform -1 0 25668 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_271
timestamp 1623529830
transform 1 0 26036 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1623529830
transform 1 0 26496 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _175_
timestamp 1623529830
transform 1 0 26128 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1623529830
transform 1 0 26220 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_279
timestamp 1623529830
transform 1 0 26772 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_283
timestamp 1623529830
transform 1 0 27140 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _136_
timestamp 1623529830
transform 1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_286
timestamp 1623529830
transform 1 0 27416 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_291
timestamp 1623529830
transform 1 0 27876 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_289
timestamp 1623529830
transform 1 0 27692 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1623529830
transform 1 0 27324 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1623529830
transform 1 0 27784 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp 1623529830
transform 1 0 27784 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_300
timestamp 1623529830
transform 1 0 28704 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_293
timestamp 1623529830
transform 1 0 28060 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_298
timestamp 1623529830
transform 1 0 28520 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _174_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform -1 0 28520 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp 1623529830
transform 1 0 28428 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform -1 0 29808 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output6
timestamp 1623529830
transform -1 0 29256 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _179_
timestamp 1623529830
transform 1 0 29624 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1623529830
transform 1 0 30452 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1623529830
transform 1 0 30176 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_306
timestamp 1623529830
transform 1 0 29256 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_313
timestamp 1623529830
transform 1 0 29900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_320
timestamp 1623529830
transform 1 0 30544 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_312
timestamp 1623529830
transform 1 0 29808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_319
timestamp 1623529830
transform 1 0 30452 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1623529830
transform 1 0 33120 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1623529830
transform 1 0 32568 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_332
timestamp 1623529830
transform 1 0 31648 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_344
timestamp 1623529830
transform 1 0 32752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1623529830
transform 1 0 33212 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_331
timestamp 1623529830
transform 1 0 31556 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_339
timestamp 1623529830
transform 1 0 32292 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_343
timestamp 1623529830
transform 1 0 32660 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output4
timestamp 1623529830
transform -1 0 33948 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_357
timestamp 1623529830
transform 1 0 33948 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_369
timestamp 1623529830
transform 1 0 35052 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_355
timestamp 1623529830
transform 1 0 33764 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_367
timestamp 1623529830
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _183_
timestamp 1623529830
transform 1 0 37076 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1623529830
transform 1 0 35788 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_378
timestamp 1623529830
transform 1 0 35880 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_390
timestamp 1623529830
transform 1 0 36984 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_379
timestamp 1623529830
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_391
timestamp 1623529830
transform 1 0 37076 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1623529830
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1623529830
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1623529830
transform 1 0 38456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1623529830
transform 1 0 37812 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output5
timestamp 1623529830
transform -1 0 38088 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_394
timestamp 1623529830
transform 1 0 37352 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_402
timestamp 1623529830
transform 1 0 38088 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_400
timestamp 1623529830
transform 1 0 37904 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_406
timestamp 1623529830
transform 1 0 38456 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1623529830
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1623529830
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1623529830
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1623529830
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_30
timestamp 1623529830
transform 1 0 3864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_42
timestamp 1623529830
transform 1 0 4968 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_54
timestamp 1623529830
transform 1 0 6072 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1623529830
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_66
timestamp 1623529830
transform 1 0 7176 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_78
timestamp 1623529830
transform 1 0 8280 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_87
timestamp 1623529830
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_99
timestamp 1623529830
transform 1 0 10212 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_111
timestamp 1623529830
transform 1 0 11316 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1623529830
transform 1 0 12420 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1623529830
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_135
timestamp 1623529830
transform 1 0 13524 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_144
timestamp 1623529830
transform 1 0 14352 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1623529830
transform -1 0 16928 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1623529830
transform 1 0 16008 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_156
timestamp 1623529830
transform 1 0 15456 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_165
timestamp 1623529830
transform 1 0 16284 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_172
timestamp 1623529830
transform 1 0 16928 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _239_
timestamp 1623529830
transform 1 0 17296 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_2_196
timestamp 1623529830
transform 1 0 19136 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _211_
timestamp 1623529830
transform -1 0 22172 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1623529830
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_201
timestamp 1623529830
transform 1 0 19596 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _205_
timestamp 1623529830
transform 1 0 22540 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_2_229
timestamp 1623529830
transform 1 0 22172 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _238_
timestamp 1623529830
transform 1 0 25208 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1623529830
transform 1 0 24748 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_253
timestamp 1623529830
transform 1 0 24380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_258
timestamp 1623529830
transform 1 0 24840 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_282
timestamp 1623529830
transform 1 0 27048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1623529830
transform -1 0 27692 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1623529830
transform 1 0 28060 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 1623529830
transform 1 0 28704 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_289
timestamp 1623529830
transform 1 0 27692 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_296
timestamp 1623529830
transform 1 0 28336 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_303
timestamp 1623529830
transform 1 0 28980 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _150_
timestamp 1623529830
transform 1 0 29348 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1623529830
transform 1 0 29992 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_310
timestamp 1623529830
transform 1 0 29624 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_315
timestamp 1623529830
transform 1 0 30084 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_327
timestamp 1623529830
transform 1 0 31188 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_339
timestamp 1623529830
transform 1 0 32292 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1623529830
transform 1 0 35236 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_351
timestamp 1623529830
transform 1 0 33396 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_363
timestamp 1623529830
transform 1 0 34500 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_372
timestamp 1623529830
transform 1 0 35328 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_384
timestamp 1623529830
transform 1 0 36432 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1623529830
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_396
timestamp 1623529830
transform 1 0 37536 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_404
timestamp 1623529830
transform 1 0 38272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1623529830
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1623529830
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1623529830
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1623529830
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1623529830
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1623529830
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_51
timestamp 1623529830
transform 1 0 5796 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_58
timestamp 1623529830
transform 1 0 6440 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_70
timestamp 1623529830
transform 1 0 7544 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_82
timestamp 1623529830
transform 1 0 8648 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_94
timestamp 1623529830
transform 1 0 9752 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_106
timestamp 1623529830
transform 1 0 10856 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1623529830
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_115
timestamp 1623529830
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_127
timestamp 1623529830
transform 1 0 12788 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_Clk
timestamp 1623529830
transform -1 0 15180 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_139
timestamp 1623529830
transform 1 0 13892 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_147
timestamp 1623529830
transform 1 0 14628 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1623529830
transform 1 0 16192 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1623529830
transform -1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1623529830
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_153
timestamp 1623529830
transform 1 0 15180 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_160
timestamp 1623529830
transform 1 0 15824 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_167
timestamp 1623529830
transform 1 0 16468 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_172
timestamp 1623529830
transform 1 0 16928 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _231_
timestamp 1623529830
transform 1 0 17664 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _208_
timestamp 1623529830
transform 1 0 19872 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_3_200
timestamp 1623529830
transform 1 0 19504 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _204_
timestamp 1623529830
transform -1 0 24472 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1623529830
transform 1 0 22080 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_224
timestamp 1623529830
transform 1 0 21712 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_229
timestamp 1623529830
transform 1 0 22172 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_233
timestamp 1623529830
transform 1 0 22540 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _200_
timestamp 1623529830
transform 1 0 24932 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_3_254
timestamp 1623529830
transform 1 0 24472 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_258
timestamp 1623529830
transform 1 0 24840 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_279
timestamp 1623529830
transform 1 0 26772 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 1623529830
transform 1 0 28888 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _177_
timestamp 1623529830
transform 1 0 27784 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1623529830
transform 1 0 27324 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_286
timestamp 1623529830
transform 1 0 27416 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_298
timestamp 1623529830
transform 1 0 28520 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_305
timestamp 1623529830
transform 1 0 29164 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _142_
timestamp 1623529830
transform 1 0 29532 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1623529830
transform 1 0 30176 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_312
timestamp 1623529830
transform 1 0 29808 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_319
timestamp 1623529830
transform 1 0 30452 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1623529830
transform 1 0 32568 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_331
timestamp 1623529830
transform 1 0 31556 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_339
timestamp 1623529830
transform 1 0 32292 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_343
timestamp 1623529830
transform 1 0 32660 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_355
timestamp 1623529830
transform 1 0 33764 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_367
timestamp 1623529830
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_379
timestamp 1623529830
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_391
timestamp 1623529830
transform 1 0 37076 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1623529830
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1623529830
transform 1 0 37812 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_400
timestamp 1623529830
transform 1 0 37904 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_406
timestamp 1623529830
transform 1 0 38456 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1623529830
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1623529830
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1623529830
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1623529830
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1623529830
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_30
timestamp 1623529830
transform 1 0 3864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_42
timestamp 1623529830
transform 1 0 4968 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_54
timestamp 1623529830
transform 1 0 6072 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1623529830
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_66
timestamp 1623529830
transform 1 0 7176 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_78
timestamp 1623529830
transform 1 0 8280 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_87
timestamp 1623529830
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_99
timestamp 1623529830
transform 1 0 10212 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_111
timestamp 1623529830
transform 1 0 11316 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1623529830
transform 1 0 12420 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _241_
timestamp 1623529830
transform -1 0 16928 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1623529830
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_135
timestamp 1623529830
transform 1 0 13524 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_144
timestamp 1623529830
transform 1 0 14352 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_172
timestamp 1623529830
transform 1 0 16928 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _229_
timestamp 1623529830
transform 1 0 17296 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_4_196
timestamp 1623529830
transform 1 0 19136 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _210_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform -1 0 21896 0 -1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1623529830
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_201
timestamp 1623529830
transform 1 0 19596 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _202_
timestamp 1623529830
transform 1 0 22540 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_4_226
timestamp 1623529830
transform 1 0 21896 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_232
timestamp 1623529830
transform 1 0 22448 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1623529830
transform 1 0 24748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_253
timestamp 1623529830
transform 1 0 24380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_258
timestamp 1623529830
transform 1 0 24840 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfstp_1  _247_
timestamp 1623529830
transform -1 0 27508 0 -1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1623529830
transform 1 0 28980 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _176_
timestamp 1623529830
transform 1 0 27876 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_287
timestamp 1623529830
transform 1 0 27508 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_299
timestamp 1623529830
transform 1 0 28612 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _144_
timestamp 1623529830
transform 1 0 30452 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1623529830
transform 1 0 29992 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_306
timestamp 1623529830
transform 1 0 29256 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_315
timestamp 1623529830
transform 1 0 30084 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_322
timestamp 1623529830
transform 1 0 30728 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_334
timestamp 1623529830
transform 1 0 31832 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_346
timestamp 1623529830
transform 1 0 32936 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1623529830
transform 1 0 35236 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_358
timestamp 1623529830
transform 1 0 34040 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_370
timestamp 1623529830
transform 1 0 35144 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_372
timestamp 1623529830
transform 1 0 35328 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_384
timestamp 1623529830
transform 1 0 36432 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1623529830
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_396
timestamp 1623529830
transform 1 0 37536 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_404
timestamp 1623529830
transform 1 0 38272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1623529830
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1623529830
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1623529830
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1623529830
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1623529830
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1623529830
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_51
timestamp 1623529830
transform 1 0 5796 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_58
timestamp 1623529830
transform 1 0 6440 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_70
timestamp 1623529830
transform 1 0 7544 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_82
timestamp 1623529830
transform 1 0 8648 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_94
timestamp 1623529830
transform 1 0 9752 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_106
timestamp 1623529830
transform 1 0 10856 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1623529830
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_115
timestamp 1623529830
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_127
timestamp 1623529830
transform 1 0 12788 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1623529830
transform -1 0 14260 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _240_
timestamp 1623529830
transform 1 0 14628 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_5_139
timestamp 1623529830
transform 1 0 13892 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_143
timestamp 1623529830
transform 1 0 14260 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1623529830
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_167
timestamp 1623529830
transform 1 0 16468 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_172
timestamp 1623529830
transform 1 0 16928 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _227_
timestamp 1623529830
transform -1 0 19504 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _206_
timestamp 1623529830
transform 1 0 19872 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_5_200
timestamp 1623529830
transform 1 0 19504 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _196_
timestamp 1623529830
transform 1 0 22632 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1623529830
transform 1 0 22080 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_224
timestamp 1623529830
transform 1 0 21712 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_229
timestamp 1623529830
transform 1 0 22172 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_233
timestamp 1623529830
transform 1 0 22540 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _199_
timestamp 1623529830
transform -1 0 26680 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_5_254
timestamp 1623529830
transform 1 0 24472 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_278
timestamp 1623529830
transform 1 0 26680 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _248_
timestamp 1623529830
transform -1 0 29624 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1623529830
transform 1 0 27324 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_284
timestamp 1623529830
transform 1 0 27232 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_286
timestamp 1623529830
transform 1 0 27416 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _135_
timestamp 1623529830
transform -1 0 30268 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _143_
timestamp 1623529830
transform 1 0 30636 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_310
timestamp 1623529830
transform 1 0 29624 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_317
timestamp 1623529830
transform 1 0 30268 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_324
timestamp 1623529830
transform 1 0 30912 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 1623529830
transform 1 0 31280 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1623529830
transform 1 0 32568 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_331
timestamp 1623529830
transform 1 0 31556 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_339
timestamp 1623529830
transform 1 0 32292 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_343
timestamp 1623529830
transform 1 0 32660 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_355
timestamp 1623529830
transform 1 0 33764 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_367
timestamp 1623529830
transform 1 0 34868 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_379
timestamp 1623529830
transform 1 0 35972 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_391
timestamp 1623529830
transform 1 0 37076 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1623529830
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1623529830
transform 1 0 37812 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_400
timestamp 1623529830
transform 1 0 37904 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_406
timestamp 1623529830
transform 1 0 38456 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1623529830
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1623529830
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1623529830
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1623529830
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1623529830
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1623529830
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1623529830
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1623529830
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_30
timestamp 1623529830
transform 1 0 3864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_42
timestamp 1623529830
transform 1 0 4968 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1623529830
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1623529830
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1623529830
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_54
timestamp 1623529830
transform 1 0 6072 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_51
timestamp 1623529830
transform 1 0 5796 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_58
timestamp 1623529830
transform 1 0 6440 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1623529830
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_66
timestamp 1623529830
transform 1 0 7176 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_78
timestamp 1623529830
transform 1 0 8280 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_87
timestamp 1623529830
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_70
timestamp 1623529830
transform 1 0 7544 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_82
timestamp 1623529830
transform 1 0 8648 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_99
timestamp 1623529830
transform 1 0 10212 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_94
timestamp 1623529830
transform 1 0 9752 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_106
timestamp 1623529830
transform 1 0 10856 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1623529830
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_111
timestamp 1623529830
transform 1 0 11316 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_123
timestamp 1623529830
transform 1 0 12420 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_115
timestamp 1623529830
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_127
timestamp 1623529830
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_139
timestamp 1623529830
transform 1 0 13892 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_139
timestamp 1623529830
transform 1 0 13892 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_135
timestamp 1623529830
transform 1 0 13524 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1623529830
transform -1 0 13892 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1623529830
transform -1 0 14260 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_143
timestamp 1623529830
transform 1 0 14260 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_144
timestamp 1623529830
transform 1 0 14352 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1623529830
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _235_
timestamp 1623529830
transform -1 0 16468 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _232_
timestamp 1623529830
transform -1 0 16928 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1623529830
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_172
timestamp 1623529830
transform 1 0 16928 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_167
timestamp 1623529830
transform 1 0 16468 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_172
timestamp 1623529830
transform 1 0 16928 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _215_
timestamp 1623529830
transform 1 0 17664 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _226_
timestamp 1623529830
transform -1 0 19136 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_6_196
timestamp 1623529830
transform 1 0 19136 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _203_
timestamp 1623529830
transform 1 0 20240 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _212_
timestamp 1623529830
transform 1 0 19872 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1623529830
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_201
timestamp 1623529830
transform 1 0 19596 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_207
timestamp 1623529830
transform 1 0 20148 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_200
timestamp 1623529830
transform 1 0 19504 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _191_
timestamp 1623529830
transform 1 0 22540 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _194_
timestamp 1623529830
transform 1 0 22448 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1623529830
transform 1 0 22080 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_228
timestamp 1623529830
transform 1 0 22080 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_224
timestamp 1623529830
transform 1 0 21712 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_229
timestamp 1623529830
transform 1 0 22172 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _197_
timestamp 1623529830
transform -1 0 26588 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _198_
timestamp 1623529830
transform 1 0 25208 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1623529830
transform 1 0 24748 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_252
timestamp 1623529830
transform 1 0 24288 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_256
timestamp 1623529830
transform 1 0 24656 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_258
timestamp 1623529830
transform 1 0 24840 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_253
timestamp 1623529830
transform 1 0 24380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_282
timestamp 1623529830
transform 1 0 27048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_277
timestamp 1623529830
transform 1 0 26588 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _201_
timestamp 1623529830
transform -1 0 29256 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _233_
timestamp 1623529830
transform 1 0 27784 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1623529830
transform 1 0 27324 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_286
timestamp 1623529830
transform 1 0 27416 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_310
timestamp 1623529830
transform 1 0 29624 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_306
timestamp 1623529830
transform 1 0 29256 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1623529830
transform 1 0 29992 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1623529830
transform 1 0 29992 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_317
timestamp 1623529830
transform 1 0 30268 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_322
timestamp 1623529830
transform 1 0 30728 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_315
timestamp 1623529830
transform 1 0 30084 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1623529830
transform 1 0 30636 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1623529830
transform 1 0 30452 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_324
timestamp 1623529830
transform 1 0 30912 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _141_
timestamp 1623529830
transform 1 0 31096 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_338
timestamp 1623529830
transform 1 0 32200 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_331
timestamp 1623529830
transform 1 0 31556 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_336
timestamp 1623529830
transform 1 0 32016 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_329
timestamp 1623529830
transform 1 0 31372 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 1623529830
transform 1 0 31924 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _145_
timestamp 1623529830
transform 1 0 31740 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1623529830
transform 1 0 31280 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1623529830
transform 1 0 32568 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 1623529830
transform 1 0 32384 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_343
timestamp 1623529830
transform 1 0 32660 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_343
timestamp 1623529830
transform 1 0 32660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1623529830
transform 1 0 35236 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_355
timestamp 1623529830
transform 1 0 33764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_367
timestamp 1623529830
transform 1 0 34868 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_355
timestamp 1623529830
transform 1 0 33764 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_367
timestamp 1623529830
transform 1 0 34868 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_372
timestamp 1623529830
transform 1 0 35328 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_384
timestamp 1623529830
transform 1 0 36432 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_379
timestamp 1623529830
transform 1 0 35972 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_391
timestamp 1623529830
transform 1 0 37076 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1623529830
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1623529830
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1623529830
transform 1 0 37812 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_396
timestamp 1623529830
transform 1 0 37536 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_404
timestamp 1623529830
transform 1 0 38272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_400
timestamp 1623529830
transform 1 0 37904 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_406
timestamp 1623529830
transform 1 0 38456 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1623529830
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1623529830
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1623529830
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1623529830
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1623529830
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_30
timestamp 1623529830
transform 1 0 3864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_42
timestamp 1623529830
transform 1 0 4968 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_54
timestamp 1623529830
transform 1 0 6072 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1623529830
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_66
timestamp 1623529830
transform 1 0 7176 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_78
timestamp 1623529830
transform 1 0 8280 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_87
timestamp 1623529830
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_99
timestamp 1623529830
transform 1 0 10212 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_111
timestamp 1623529830
transform 1 0 11316 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1623529830
transform 1 0 12420 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _234_
timestamp 1623529830
transform 1 0 15088 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1623529830
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_135
timestamp 1623529830
transform 1 0 13524 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_144
timestamp 1623529830
transform 1 0 14352 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_172
timestamp 1623529830
transform 1 0 16928 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _218_
timestamp 1623529830
transform 1 0 17296 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_8_196
timestamp 1623529830
transform 1 0 19136 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _213_
timestamp 1623529830
transform -1 0 21988 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1623529830
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_201
timestamp 1623529830
transform 1 0 19596 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _189_
timestamp 1623529830
transform -1 0 24196 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_8_227
timestamp 1623529830
transform 1 0 21988 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _195_
timestamp 1623529830
transform -1 0 27048 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1623529830
transform 1 0 24748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_251
timestamp 1623529830
transform 1 0 24196 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_258
timestamp 1623529830
transform 1 0 24840 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_282
timestamp 1623529830
transform 1 0 27048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _222_
timestamp 1623529830
transform 1 0 27416 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1623529830
transform 1 0 30452 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _147_
timestamp 1623529830
transform 1 0 31096 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1623529830
transform 1 0 29992 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_306
timestamp 1623529830
transform 1 0 29256 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_315
timestamp 1623529830
transform 1 0 30084 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_322
timestamp 1623529830
transform 1 0 30728 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1623529830
transform 1 0 31740 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_Clk
timestamp 1623529830
transform 1 0 32384 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_329
timestamp 1623529830
transform 1 0 31372 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_336
timestamp 1623529830
transform 1 0 32016 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_343
timestamp 1623529830
transform 1 0 32660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1623529830
transform 1 0 35236 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_355
timestamp 1623529830
transform 1 0 33764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_367
timestamp 1623529830
transform 1 0 34868 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_372
timestamp 1623529830
transform 1 0 35328 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_384
timestamp 1623529830
transform 1 0 36432 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1623529830
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_396
timestamp 1623529830
transform 1 0 37536 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_404
timestamp 1623529830
transform 1 0 38272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1623529830
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1623529830
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1623529830
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1623529830
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1623529830
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1623529830
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_51
timestamp 1623529830
transform 1 0 5796 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_58
timestamp 1623529830
transform 1 0 6440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_70
timestamp 1623529830
transform 1 0 7544 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_82
timestamp 1623529830
transform 1 0 8648 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_94
timestamp 1623529830
transform 1 0 9752 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_106
timestamp 1623529830
transform 1 0 10856 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1623529830
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_115
timestamp 1623529830
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_127
timestamp 1623529830
transform 1 0 12788 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_Clk
timestamp 1623529830
transform -1 0 15180 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_139
timestamp 1623529830
transform 1 0 13892 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_147
timestamp 1623529830
transform 1 0 14628 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1623529830
transform -1 0 16468 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1623529830
transform -1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1623529830
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_153
timestamp 1623529830
transform 1 0 15180 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_160
timestamp 1623529830
transform 1 0 15824 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_167
timestamp 1623529830
transform 1 0 16468 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_172
timestamp 1623529830
transform 1 0 16928 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _221_
timestamp 1623529830
transform 1 0 17664 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _214_
timestamp 1623529830
transform 1 0 19872 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_9_200
timestamp 1623529830
transform 1 0 19504 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _187_
timestamp 1623529830
transform -1 0 24564 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1623529830
transform 1 0 22080 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_224
timestamp 1623529830
transform 1 0 21712 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_229
timestamp 1623529830
transform 1 0 22172 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _193_
timestamp 1623529830
transform -1 0 26772 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_9_255
timestamp 1623529830
transform 1 0 24564 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_279
timestamp 1623529830
transform 1 0 26772 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _249_
timestamp 1623529830
transform 1 0 27784 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1623529830
transform 1 0 27324 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_286
timestamp 1623529830
transform 1 0 27416 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _129_
timestamp 1623529830
transform 1 0 29992 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _152_
timestamp 1623529830
transform 1 0 30636 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_310
timestamp 1623529830
transform 1 0 29624 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_317
timestamp 1623529830
transform 1 0 30268 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_324
timestamp 1623529830
transform 1 0 30912 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1623529830
transform 1 0 31280 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1623529830
transform 1 0 32568 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_331
timestamp 1623529830
transform 1 0 31556 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_339
timestamp 1623529830
transform 1 0 32292 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_343
timestamp 1623529830
transform 1 0 32660 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_355
timestamp 1623529830
transform 1 0 33764 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_367
timestamp 1623529830
transform 1 0 34868 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_379
timestamp 1623529830
transform 1 0 35972 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_391
timestamp 1623529830
transform 1 0 37076 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1623529830
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1623529830
transform 1 0 37812 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_400
timestamp 1623529830
transform 1 0 37904 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_406
timestamp 1623529830
transform 1 0 38456 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1623529830
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1623529830
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1623529830
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1623529830
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1623529830
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1623529830
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1623529830
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_54
timestamp 1623529830
transform 1 0 6072 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1623529830
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_66
timestamp 1623529830
transform 1 0 7176 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_78
timestamp 1623529830
transform 1 0 8280 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_87
timestamp 1623529830
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_99
timestamp 1623529830
transform 1 0 10212 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_111
timestamp 1623529830
transform 1 0 11316 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1623529830
transform 1 0 12420 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1623529830
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_135
timestamp 1623529830
transform 1 0 13524 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_144
timestamp 1623529830
transform 1 0 14352 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1623529830
transform 1 0 16652 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_Clk
timestamp 1623529830
transform -1 0 16284 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_156
timestamp 1623529830
transform 1 0 15456 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_165
timestamp 1623529830
transform 1 0 16284 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_172
timestamp 1623529830
transform 1 0 16928 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _224_
timestamp 1623529830
transform 1 0 17296 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_10_196
timestamp 1623529830
transform 1 0 19136 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _192_
timestamp 1623529830
transform 1 0 20332 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1623529830
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_201
timestamp 1623529830
transform 1 0 19596 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _186_
timestamp 1623529830
transform 1 0 22540 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_10_229
timestamp 1623529830
transform 1 0 22172 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _217_
timestamp 1623529830
transform 1 0 25208 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1623529830
transform 1 0 24748 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_253
timestamp 1623529830
transform 1 0 24380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_258
timestamp 1623529830
transform 1 0 24840 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_282
timestamp 1623529830
transform 1 0 27048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _252_
timestamp 1623529830
transform -1 0 29256 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1623529830
transform 1 0 30452 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1623529830
transform 1 0 29992 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_Clk
timestamp 1623529830
transform 1 0 31096 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_306
timestamp 1623529830
transform 1 0 29256 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_315
timestamp 1623529830
transform 1 0 30084 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_322
timestamp 1623529830
transform 1 0 30728 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_329
timestamp 1623529830
transform 1 0 31372 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_341
timestamp 1623529830
transform 1 0 32476 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1623529830
transform 1 0 35236 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_353
timestamp 1623529830
transform 1 0 33580 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_365
timestamp 1623529830
transform 1 0 34684 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_372
timestamp 1623529830
transform 1 0 35328 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_384
timestamp 1623529830
transform 1 0 36432 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1623529830
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_396
timestamp 1623529830
transform 1 0 37536 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_404
timestamp 1623529830
transform 1 0 38272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1623529830
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1623529830
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1623529830
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1623529830
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1623529830
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1623529830
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_51
timestamp 1623529830
transform 1 0 5796 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_58
timestamp 1623529830
transform 1 0 6440 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_70
timestamp 1623529830
transform 1 0 7544 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_82
timestamp 1623529830
transform 1 0 8648 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_94
timestamp 1623529830
transform 1 0 9752 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_106
timestamp 1623529830
transform 1 0 10856 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1623529830
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_115
timestamp 1623529830
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_127
timestamp 1623529830
transform 1 0 12788 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_139
timestamp 1623529830
transform 1 0 13892 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_151
timestamp 1623529830
transform 1 0 14996 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1623529830
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_163
timestamp 1623529830
transform 1 0 16100 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_172
timestamp 1623529830
transform 1 0 16928 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _225_
timestamp 1623529830
transform -1 0 19504 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _216_
timestamp 1623529830
transform -1 0 21712 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_11_200
timestamp 1623529830
transform 1 0 19504 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _185_
timestamp 1623529830
transform 1 0 23000 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1623529830
transform 1 0 22080 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_224
timestamp 1623529830
transform 1 0 21712 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_229
timestamp 1623529830
transform 1 0 22172 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_237
timestamp 1623529830
transform 1 0 22908 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _092_
timestamp 1623529830
transform 1 0 25208 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_258
timestamp 1623529830
transform 1 0 24840 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1623529830
transform 1 0 25852 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1623529830
transform 1 0 26496 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_265
timestamp 1623529830
transform 1 0 25484 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_272
timestamp 1623529830
transform 1 0 26128 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_279
timestamp 1623529830
transform 1 0 26772 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _253_
timestamp 1623529830
transform 1 0 27784 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1623529830
transform 1 0 27324 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_286
timestamp 1623529830
transform 1 0 27416 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1623529830
transform 1 0 29992 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_310
timestamp 1623529830
transform 1 0 29624 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1623529830
transform 1 0 30268 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1623529830
transform 1 0 32568 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_329
timestamp 1623529830
transform 1 0 31372 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_341
timestamp 1623529830
transform 1 0 32476 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_343
timestamp 1623529830
transform 1 0 32660 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_355
timestamp 1623529830
transform 1 0 33764 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_367
timestamp 1623529830
transform 1 0 34868 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_379
timestamp 1623529830
transform 1 0 35972 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_391
timestamp 1623529830
transform 1 0 37076 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1623529830
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1623529830
transform 1 0 37812 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_400
timestamp 1623529830
transform 1 0 37904 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_406
timestamp 1623529830
transform 1 0 38456 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1623529830
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1623529830
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1623529830
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1623529830
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1623529830
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_30
timestamp 1623529830
transform 1 0 3864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_42
timestamp 1623529830
transform 1 0 4968 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_54
timestamp 1623529830
transform 1 0 6072 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1623529830
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_66
timestamp 1623529830
transform 1 0 7176 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_78
timestamp 1623529830
transform 1 0 8280 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_87
timestamp 1623529830
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_99
timestamp 1623529830
transform 1 0 10212 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_111
timestamp 1623529830
transform 1 0 11316 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_123
timestamp 1623529830
transform 1 0 12420 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1623529830
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_135
timestamp 1623529830
transform 1 0 13524 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_144
timestamp 1623529830
transform 1 0 14352 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_156
timestamp 1623529830
transform 1 0 15456 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_168
timestamp 1623529830
transform 1 0 16560 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1623529830
transform -1 0 19136 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1623529830
transform -1 0 18492 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _122_
timestamp 1623529830
transform 1 0 17572 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_176
timestamp 1623529830
transform 1 0 17296 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_182
timestamp 1623529830
transform 1 0 17848 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_189
timestamp 1623529830
transform 1 0 18492 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_196
timestamp 1623529830
transform 1 0 19136 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _220_
timestamp 1623529830
transform 1 0 20240 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1623529830
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_201
timestamp 1623529830
transform 1 0 19596 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_207
timestamp 1623529830
transform 1 0 20148 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _188_
timestamp 1623529830
transform 1 0 22448 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_12_228
timestamp 1623529830
transform 1 0 22080 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _250_
timestamp 1623529830
transform 1 0 25208 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1623529830
transform 1 0 24748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_252
timestamp 1623529830
transform 1 0 24288 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_256
timestamp 1623529830
transform 1 0 24656 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_258
timestamp 1623529830
transform 1 0 24840 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_282
timestamp 1623529830
transform 1 0 27048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1623529830
transform 1 0 27416 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1623529830
transform 1 0 28060 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1623529830
transform 1 0 28704 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_289
timestamp 1623529830
transform 1 0 27692 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_296
timestamp 1623529830
transform 1 0 28336 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_303
timestamp 1623529830
transform 1 0 28980 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1623529830
transform 1 0 29992 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_311
timestamp 1623529830
transform 1 0 29716 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_315
timestamp 1623529830
transform 1 0 30084 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_327
timestamp 1623529830
transform 1 0 31188 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_339
timestamp 1623529830
transform 1 0 32292 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1623529830
transform 1 0 35236 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_351
timestamp 1623529830
transform 1 0 33396 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_363
timestamp 1623529830
transform 1 0 34500 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_372
timestamp 1623529830
transform 1 0 35328 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_384
timestamp 1623529830
transform 1 0 36432 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1623529830
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_396
timestamp 1623529830
transform 1 0 37536 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_404
timestamp 1623529830
transform 1 0 38272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1623529830
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1623529830
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1623529830
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1623529830
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1623529830
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1623529830
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1623529830
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1623529830
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1623529830
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1623529830
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1623529830
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_42
timestamp 1623529830
transform 1 0 4968 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1623529830
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_51
timestamp 1623529830
transform 1 0 5796 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_58
timestamp 1623529830
transform 1 0 6440 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_54
timestamp 1623529830
transform 1 0 6072 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1623529830
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_70
timestamp 1623529830
transform 1 0 7544 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_82
timestamp 1623529830
transform 1 0 8648 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_66
timestamp 1623529830
transform 1 0 7176 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_78
timestamp 1623529830
transform 1 0 8280 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_87
timestamp 1623529830
transform 1 0 9108 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_94
timestamp 1623529830
transform 1 0 9752 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_106
timestamp 1623529830
transform 1 0 10856 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_99
timestamp 1623529830
transform 1 0 10212 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1623529830
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_115
timestamp 1623529830
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_127
timestamp 1623529830
transform 1 0 12788 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_111
timestamp 1623529830
transform 1 0 11316 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_123
timestamp 1623529830
transform 1 0 12420 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1623529830
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_139
timestamp 1623529830
transform 1 0 13892 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_151
timestamp 1623529830
transform 1 0 14996 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_135
timestamp 1623529830
transform 1 0 13524 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_144
timestamp 1623529830
transform 1 0 14352 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1623529830
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_163
timestamp 1623529830
transform 1 0 16100 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_172
timestamp 1623529830
transform 1 0 16928 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_156
timestamp 1623529830
transform 1 0 15456 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_168
timestamp 1623529830
transform 1 0 16560 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1623529830
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_Clk
timestamp 1623529830
transform 1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_184
timestamp 1623529830
transform 1 0 18032 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_193
timestamp 1623529830
transform 1 0 18860 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_180
timestamp 1623529830
transform 1 0 17664 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_192
timestamp 1623529830
transform 1 0 18768 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_196
timestamp 1623529830
transform 1 0 19136 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _097_
timestamp 1623529830
transform -1 0 21068 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1623529830
transform 1 0 20148 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1623529830
transform -1 0 19504 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _223_
timestamp 1623529830
transform 1 0 19872 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1623529830
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_200
timestamp 1623529830
transform 1 0 19504 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_201
timestamp 1623529830
transform 1 0 19596 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_210
timestamp 1623529830
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_217
timestamp 1623529830
transform 1 0 21068 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _190_
timestamp 1623529830
transform 1 0 22540 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _219_
timestamp 1623529830
transform -1 0 23276 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1623529830
transform 1 0 22080 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_224
timestamp 1623529830
transform 1 0 21712 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_229
timestamp 1623529830
transform 1 0 22172 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _091_
timestamp 1623529830
transform 1 0 23644 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1623529830
transform 1 0 25208 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _251_
timestamp 1623529830
transform -1 0 26588 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1623529830
transform 1 0 24748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_253
timestamp 1623529830
transform 1 0 24380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_241
timestamp 1623529830
transform 1 0 23276 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_248
timestamp 1623529830
transform 1 0 23920 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_256
timestamp 1623529830
transform 1 0 24656 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_258
timestamp 1623529830
transform 1 0 24840 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1623529830
transform 1 0 25852 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _157_
timestamp 1623529830
transform 1 0 26496 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1623529830
transform 1 0 27140 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_277
timestamp 1623529830
transform 1 0 26588 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_265
timestamp 1623529830
transform 1 0 25484 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_272
timestamp 1623529830
transform 1 0 26128 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_279
timestamp 1623529830
transform 1 0 26772 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_286
timestamp 1623529830
transform 1 0 27416 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_293
timestamp 1623529830
transform 1 0 28060 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_286
timestamp 1623529830
transform 1 0 27416 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_Clk
timestamp 1623529830
transform -1 0 28060 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1623529830
transform 1 0 27324 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1623529830
transform 1 0 27784 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_305
timestamp 1623529830
transform 1 0 29164 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1623529830
transform 1 0 28428 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_293
timestamp 1623529830
transform 1 0 28060 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_300
timestamp 1623529830
transform 1 0 28704 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1623529830
transform 1 0 29992 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_312
timestamp 1623529830
transform 1 0 29808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_324
timestamp 1623529830
transform 1 0 30912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_313
timestamp 1623529830
transform 1 0 29900 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_315
timestamp 1623529830
transform 1 0 30084 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_327
timestamp 1623529830
transform 1 0 31188 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1623529830
transform 1 0 32568 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_336
timestamp 1623529830
transform 1 0 32016 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_343
timestamp 1623529830
transform 1 0 32660 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_339
timestamp 1623529830
transform 1 0 32292 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1623529830
transform 1 0 35236 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_355
timestamp 1623529830
transform 1 0 33764 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_367
timestamp 1623529830
transform 1 0 34868 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_351
timestamp 1623529830
transform 1 0 33396 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_363
timestamp 1623529830
transform 1 0 34500 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_379
timestamp 1623529830
transform 1 0 35972 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_391
timestamp 1623529830
transform 1 0 37076 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_372
timestamp 1623529830
transform 1 0 35328 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_384
timestamp 1623529830
transform 1 0 36432 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1623529830
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1623529830
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1623529830
transform 1 0 37812 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_400
timestamp 1623529830
transform 1 0 37904 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_406
timestamp 1623529830
transform 1 0 38456 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_396
timestamp 1623529830
transform 1 0 37536 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_404
timestamp 1623529830
transform 1 0 38272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1623529830
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1623529830
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1623529830
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1623529830
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1623529830
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1623529830
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_51
timestamp 1623529830
transform 1 0 5796 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_58
timestamp 1623529830
transform 1 0 6440 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_70
timestamp 1623529830
transform 1 0 7544 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_82
timestamp 1623529830
transform 1 0 8648 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_94
timestamp 1623529830
transform 1 0 9752 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_106
timestamp 1623529830
transform 1 0 10856 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1623529830
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_115
timestamp 1623529830
transform 1 0 11684 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_127
timestamp 1623529830
transform 1 0 12788 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_139
timestamp 1623529830
transform 1 0 13892 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_151
timestamp 1623529830
transform 1 0 14996 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1623529830
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_163
timestamp 1623529830
transform 1 0 16100 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_172
timestamp 1623529830
transform 1 0 16928 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_Clk
timestamp 1623529830
transform 1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_184
timestamp 1623529830
transform 1 0 18032 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_192
timestamp 1623529830
transform 1 0 18768 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1623529830
transform 1 0 19136 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _110_
timestamp 1623529830
transform -1 0 21068 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1623529830
transform 1 0 20148 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_Clk
timestamp 1623529830
transform 1 0 19504 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_203
timestamp 1623529830
transform 1 0 19780 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_210
timestamp 1623529830
transform 1 0 20424 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_217
timestamp 1623529830
transform 1 0 21068 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _104_
timestamp 1623529830
transform -1 0 21712 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _237_
timestamp 1623529830
transform -1 0 24380 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1623529830
transform 1 0 22080 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_224
timestamp 1623529830
transform 1 0 21712 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_229
timestamp 1623529830
transform 1 0 22172 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1623529830
transform 1 0 24748 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_253
timestamp 1623529830
transform 1 0 24380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_260
timestamp 1623529830
transform 1 0 25024 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _128_
timestamp 1623529830
transform 1 0 25392 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1623529830
transform 1 0 26036 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_267
timestamp 1623529830
transform 1 0 25668 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_274
timestamp 1623529830
transform 1 0 26312 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_282
timestamp 1623529830
transform 1 0 27048 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1623529830
transform 1 0 27324 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_286
timestamp 1623529830
transform 1 0 27416 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_298
timestamp 1623529830
transform 1 0 28520 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_310
timestamp 1623529830
transform 1 0 29624 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_322
timestamp 1623529830
transform 1 0 30728 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1623529830
transform 1 0 32568 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_334
timestamp 1623529830
transform 1 0 31832 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_343
timestamp 1623529830
transform 1 0 32660 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_355
timestamp 1623529830
transform 1 0 33764 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_367
timestamp 1623529830
transform 1 0 34868 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_379
timestamp 1623529830
transform 1 0 35972 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_391
timestamp 1623529830
transform 1 0 37076 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1623529830
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1623529830
transform 1 0 37812 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_400
timestamp 1623529830
transform 1 0 37904 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_406
timestamp 1623529830
transform 1 0 38456 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1623529830
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1623529830
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1623529830
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1623529830
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1623529830
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_30
timestamp 1623529830
transform 1 0 3864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_42
timestamp 1623529830
transform 1 0 4968 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_54
timestamp 1623529830
transform 1 0 6072 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1623529830
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_66
timestamp 1623529830
transform 1 0 7176 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_78
timestamp 1623529830
transform 1 0 8280 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_87
timestamp 1623529830
transform 1 0 9108 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_99
timestamp 1623529830
transform 1 0 10212 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_111
timestamp 1623529830
transform 1 0 11316 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_123
timestamp 1623529830
transform 1 0 12420 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1623529830
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_135
timestamp 1623529830
transform 1 0 13524 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_144
timestamp 1623529830
transform 1 0 14352 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_156
timestamp 1623529830
transform 1 0 15456 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_168
timestamp 1623529830
transform 1 0 16560 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_180
timestamp 1623529830
transform 1 0 17664 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_192
timestamp 1623529830
transform 1 0 18768 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _236_
timestamp 1623529830
transform -1 0 23000 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1623529830
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_Clk
timestamp 1623529830
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_201
timestamp 1623529830
transform 1 0 19596 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_209
timestamp 1623529830
transform 1 0 20332 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_214
timestamp 1623529830
transform 1 0 20792 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_238
timestamp 1623529830
transform 1 0 23000 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1623529830
transform 1 0 23368 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1623529830
transform 1 0 24012 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _156_
timestamp 1623529830
transform -1 0 25484 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1623529830
transform 1 0 24748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_245
timestamp 1623529830
transform 1 0 23644 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_252
timestamp 1623529830
transform 1 0 24288 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_256
timestamp 1623529830
transform 1 0 24656 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_258
timestamp 1623529830
transform 1 0 24840 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_Clk
timestamp 1623529830
transform -1 0 26128 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_265
timestamp 1623529830
transform 1 0 25484 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_272
timestamp 1623529830
transform 1 0 26128 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_284
timestamp 1623529830
transform 1 0 27232 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_296
timestamp 1623529830
transform 1 0 28336 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1623529830
transform 1 0 29992 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_308
timestamp 1623529830
transform 1 0 29440 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_315
timestamp 1623529830
transform 1 0 30084 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_327
timestamp 1623529830
transform 1 0 31188 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_339
timestamp 1623529830
transform 1 0 32292 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1623529830
transform 1 0 35236 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_351
timestamp 1623529830
transform 1 0 33396 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_363
timestamp 1623529830
transform 1 0 34500 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_372
timestamp 1623529830
transform 1 0 35328 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_384
timestamp 1623529830
transform 1 0 36432 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1623529830
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_396
timestamp 1623529830
transform 1 0 37536 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_404
timestamp 1623529830
transform 1 0 38272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1623529830
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1623529830
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1623529830
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1623529830
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1623529830
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1623529830
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_51
timestamp 1623529830
transform 1 0 5796 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_58
timestamp 1623529830
transform 1 0 6440 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_70
timestamp 1623529830
transform 1 0 7544 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_82
timestamp 1623529830
transform 1 0 8648 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_94
timestamp 1623529830
transform 1 0 9752 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_106
timestamp 1623529830
transform 1 0 10856 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1623529830
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_115
timestamp 1623529830
transform 1 0 11684 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_127
timestamp 1623529830
transform 1 0 12788 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_139
timestamp 1623529830
transform 1 0 13892 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_151
timestamp 1623529830
transform 1 0 14996 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1623529830
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_163
timestamp 1623529830
transform 1 0 16100 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_172
timestamp 1623529830
transform 1 0 16928 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1623529830
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1623529830
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1623529830
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _116_
timestamp 1623529830
transform -1 0 22816 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1623529830
transform 1 0 23184 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1623529830
transform 1 0 22080 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_Clk
timestamp 1623529830
transform -1 0 21712 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_220
timestamp 1623529830
transform 1 0 21344 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_224
timestamp 1623529830
transform 1 0 21712 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_229
timestamp 1623529830
transform 1 0 22172 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_236
timestamp 1623529830
transform 1 0 22816 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _153_
timestamp 1623529830
transform 1 0 23828 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1623529830
transform 1 0 24472 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1623529830
transform 1 0 25116 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_243
timestamp 1623529830
transform 1 0 23460 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_250
timestamp 1623529830
transform 1 0 24104 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_257
timestamp 1623529830
transform 1 0 24748 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_264
timestamp 1623529830
transform 1 0 25392 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_276
timestamp 1623529830
transform 1 0 26496 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1623529830
transform 1 0 27324 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_284
timestamp 1623529830
transform 1 0 27232 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_286
timestamp 1623529830
transform 1 0 27416 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_298
timestamp 1623529830
transform 1 0 28520 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_310
timestamp 1623529830
transform 1 0 29624 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_322
timestamp 1623529830
transform 1 0 30728 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1623529830
transform 1 0 32568 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_334
timestamp 1623529830
transform 1 0 31832 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_343
timestamp 1623529830
transform 1 0 32660 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_355
timestamp 1623529830
transform 1 0 33764 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_367
timestamp 1623529830
transform 1 0 34868 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_379
timestamp 1623529830
transform 1 0 35972 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_391
timestamp 1623529830
transform 1 0 37076 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1623529830
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1623529830
transform 1 0 37812 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_400
timestamp 1623529830
transform 1 0 37904 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_406
timestamp 1623529830
transform 1 0 38456 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1623529830
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1623529830
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1623529830
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1623529830
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1623529830
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_30
timestamp 1623529830
transform 1 0 3864 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_42
timestamp 1623529830
transform 1 0 4968 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_54
timestamp 1623529830
transform 1 0 6072 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1623529830
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_66
timestamp 1623529830
transform 1 0 7176 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_78
timestamp 1623529830
transform 1 0 8280 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_87
timestamp 1623529830
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_99
timestamp 1623529830
transform 1 0 10212 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_111
timestamp 1623529830
transform 1 0 11316 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_123
timestamp 1623529830
transform 1 0 12420 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1623529830
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_135
timestamp 1623529830
transform 1 0 13524 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_144
timestamp 1623529830
transform 1 0 14352 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_156
timestamp 1623529830
transform 1 0 15456 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_168
timestamp 1623529830
transform 1 0 16560 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_180
timestamp 1623529830
transform 1 0 17664 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_192
timestamp 1623529830
transform 1 0 18768 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1623529830
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_Clk
timestamp 1623529830
transform 1 0 19964 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_201
timestamp 1623529830
transform 1 0 19596 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_208
timestamp 1623529830
transform 1 0 20240 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_Clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 21896 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_18_220
timestamp 1623529830
transform 1 0 21344 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _159_
timestamp 1623529830
transform 1 0 24104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _163_
timestamp 1623529830
transform 1 0 25208 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1623529830
transform 1 0 24748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_246
timestamp 1623529830
transform 1 0 23736 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_253
timestamp 1623529830
transform 1 0 24380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_258
timestamp 1623529830
transform 1 0 24840 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1623529830
transform 1 0 25484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1623529830
transform 1 0 26588 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1623529830
transform 1 0 27692 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_301
timestamp 1623529830
transform 1 0 28796 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1623529830
transform 1 0 29992 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_313
timestamp 1623529830
transform 1 0 29900 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_315
timestamp 1623529830
transform 1 0 30084 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_327
timestamp 1623529830
transform 1 0 31188 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_339
timestamp 1623529830
transform 1 0 32292 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1623529830
transform 1 0 35236 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_351
timestamp 1623529830
transform 1 0 33396 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_363
timestamp 1623529830
transform 1 0 34500 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_372
timestamp 1623529830
transform 1 0 35328 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_384
timestamp 1623529830
transform 1 0 36432 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1623529830
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_396
timestamp 1623529830
transform 1 0 37536 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_404
timestamp 1623529830
transform 1 0 38272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1623529830
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1623529830
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1623529830
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1623529830
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1623529830
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1623529830
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1623529830
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1623529830
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1623529830
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1623529830
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_30
timestamp 1623529830
transform 1 0 3864 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_42
timestamp 1623529830
transform 1 0 4968 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1623529830
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_51
timestamp 1623529830
transform 1 0 5796 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_58
timestamp 1623529830
transform 1 0 6440 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_54
timestamp 1623529830
transform 1 0 6072 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1623529830
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_70
timestamp 1623529830
transform 1 0 7544 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_82
timestamp 1623529830
transform 1 0 8648 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_66
timestamp 1623529830
transform 1 0 7176 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_78
timestamp 1623529830
transform 1 0 8280 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_87
timestamp 1623529830
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_94
timestamp 1623529830
transform 1 0 9752 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_106
timestamp 1623529830
transform 1 0 10856 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_99
timestamp 1623529830
transform 1 0 10212 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1623529830
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_115
timestamp 1623529830
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_127
timestamp 1623529830
transform 1 0 12788 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_111
timestamp 1623529830
transform 1 0 11316 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_123
timestamp 1623529830
transform 1 0 12420 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1623529830
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_139
timestamp 1623529830
transform 1 0 13892 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_151
timestamp 1623529830
transform 1 0 14996 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_135
timestamp 1623529830
transform 1 0 13524 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_144
timestamp 1623529830
transform 1 0 14352 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1623529830
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_163
timestamp 1623529830
transform 1 0 16100 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_172
timestamp 1623529830
transform 1 0 16928 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_156
timestamp 1623529830
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_168
timestamp 1623529830
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1623529830
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1623529830
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_180
timestamp 1623529830
transform 1 0 17664 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_192
timestamp 1623529830
transform 1 0 18768 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1623529830
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1623529830
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_201
timestamp 1623529830
transform 1 0 19596 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_213
timestamp 1623529830
transform 1 0 20700 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1623529830
transform 1 0 22080 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_220
timestamp 1623529830
transform 1 0 21344 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_229
timestamp 1623529830
transform 1 0 22172 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_225
timestamp 1623529830
transform 1 0 21804 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_237
timestamp 1623529830
transform 1 0 22908 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1623529830
transform 1 0 24748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_241
timestamp 1623529830
transform 1 0 23276 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_253
timestamp 1623529830
transform 1 0 24380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_249
timestamp 1623529830
transform 1 0 24012 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_258
timestamp 1623529830
transform 1 0 24840 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_265
timestamp 1623529830
transform 1 0 25484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_277
timestamp 1623529830
transform 1 0 26588 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_270
timestamp 1623529830
transform 1 0 25944 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_282
timestamp 1623529830
transform 1 0 27048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1623529830
transform 1 0 27324 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_286
timestamp 1623529830
transform 1 0 27416 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_298
timestamp 1623529830
transform 1 0 28520 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_294
timestamp 1623529830
transform 1 0 28152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1623529830
transform 1 0 29992 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_310
timestamp 1623529830
transform 1 0 29624 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_322
timestamp 1623529830
transform 1 0 30728 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_306
timestamp 1623529830
transform 1 0 29256 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_315
timestamp 1623529830
transform 1 0 30084 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_327
timestamp 1623529830
transform 1 0 31188 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1623529830
transform 1 0 32568 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_334
timestamp 1623529830
transform 1 0 31832 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_343
timestamp 1623529830
transform 1 0 32660 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_339
timestamp 1623529830
transform 1 0 32292 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1623529830
transform 1 0 35236 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_355
timestamp 1623529830
transform 1 0 33764 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_367
timestamp 1623529830
transform 1 0 34868 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_351
timestamp 1623529830
transform 1 0 33396 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_363
timestamp 1623529830
transform 1 0 34500 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_379
timestamp 1623529830
transform 1 0 35972 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_391
timestamp 1623529830
transform 1 0 37076 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_372
timestamp 1623529830
transform 1 0 35328 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_384
timestamp 1623529830
transform 1 0 36432 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1623529830
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1623529830
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1623529830
transform 1 0 37812 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_400
timestamp 1623529830
transform 1 0 37904 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_406
timestamp 1623529830
transform 1 0 38456 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_396
timestamp 1623529830
transform 1 0 37536 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_404
timestamp 1623529830
transform 1 0 38272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1623529830
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1623529830
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1623529830
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1623529830
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1623529830
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1623529830
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_51
timestamp 1623529830
transform 1 0 5796 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_58
timestamp 1623529830
transform 1 0 6440 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_70
timestamp 1623529830
transform 1 0 7544 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_82
timestamp 1623529830
transform 1 0 8648 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_94
timestamp 1623529830
transform 1 0 9752 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_106
timestamp 1623529830
transform 1 0 10856 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1623529830
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_115
timestamp 1623529830
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_127
timestamp 1623529830
transform 1 0 12788 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_139
timestamp 1623529830
transform 1 0 13892 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_151
timestamp 1623529830
transform 1 0 14996 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1623529830
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_163
timestamp 1623529830
transform 1 0 16100 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_172
timestamp 1623529830
transform 1 0 16928 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1623529830
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1623529830
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1623529830
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1623529830
transform 1 0 22080 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_220
timestamp 1623529830
transform 1 0 21344 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_229
timestamp 1623529830
transform 1 0 22172 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_241
timestamp 1623529830
transform 1 0 23276 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_253
timestamp 1623529830
transform 1 0 24380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_265
timestamp 1623529830
transform 1 0 25484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_277
timestamp 1623529830
transform 1 0 26588 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1623529830
transform 1 0 27324 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_286
timestamp 1623529830
transform 1 0 27416 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_298
timestamp 1623529830
transform 1 0 28520 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_310
timestamp 1623529830
transform 1 0 29624 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_322
timestamp 1623529830
transform 1 0 30728 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1623529830
transform 1 0 32568 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_334
timestamp 1623529830
transform 1 0 31832 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_343
timestamp 1623529830
transform 1 0 32660 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_355
timestamp 1623529830
transform 1 0 33764 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_367
timestamp 1623529830
transform 1 0 34868 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_379
timestamp 1623529830
transform 1 0 35972 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_391
timestamp 1623529830
transform 1 0 37076 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1623529830
transform -1 0 38824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1623529830
transform 1 0 37812 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_400
timestamp 1623529830
transform 1 0 37904 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_406
timestamp 1623529830
transform 1 0 38456 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1623529830
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1623529830
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1623529830
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1623529830
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1623529830
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_30
timestamp 1623529830
transform 1 0 3864 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_42
timestamp 1623529830
transform 1 0 4968 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_54
timestamp 1623529830
transform 1 0 6072 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1623529830
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_66
timestamp 1623529830
transform 1 0 7176 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_78
timestamp 1623529830
transform 1 0 8280 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_87
timestamp 1623529830
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_99
timestamp 1623529830
transform 1 0 10212 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_111
timestamp 1623529830
transform 1 0 11316 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_123
timestamp 1623529830
transform 1 0 12420 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1623529830
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_135
timestamp 1623529830
transform 1 0 13524 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_144
timestamp 1623529830
transform 1 0 14352 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_156
timestamp 1623529830
transform 1 0 15456 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_168
timestamp 1623529830
transform 1 0 16560 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_180
timestamp 1623529830
transform 1 0 17664 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_192
timestamp 1623529830
transform 1 0 18768 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1623529830
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_201
timestamp 1623529830
transform 1 0 19596 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_213
timestamp 1623529830
transform 1 0 20700 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _090_
timestamp 1623529830
transform 1 0 22724 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_225
timestamp 1623529830
transform 1 0 21804 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_233
timestamp 1623529830
transform 1 0 22540 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_238
timestamp 1623529830
transform 1 0 23000 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1623529830
transform 1 0 24748 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_250
timestamp 1623529830
transform 1 0 24104 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_256
timestamp 1623529830
transform 1 0 24656 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_258
timestamp 1623529830
transform 1 0 24840 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_270
timestamp 1623529830
transform 1 0 25944 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_282
timestamp 1623529830
transform 1 0 27048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_294
timestamp 1623529830
transform 1 0 28152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1623529830
transform 1 0 29992 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_306
timestamp 1623529830
transform 1 0 29256 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_315
timestamp 1623529830
transform 1 0 30084 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_327
timestamp 1623529830
transform 1 0 31188 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_339
timestamp 1623529830
transform 1 0 32292 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1623529830
transform 1 0 35236 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_351
timestamp 1623529830
transform 1 0 33396 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_363
timestamp 1623529830
transform 1 0 34500 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_372
timestamp 1623529830
transform 1 0 35328 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_384
timestamp 1623529830
transform 1 0 36432 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1623529830
transform -1 0 38824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_396
timestamp 1623529830
transform 1 0 37536 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_404
timestamp 1623529830
transform 1 0 38272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1623529830
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1623529830
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1623529830
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1623529830
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1623529830
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1623529830
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_51
timestamp 1623529830
transform 1 0 5796 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_58
timestamp 1623529830
transform 1 0 6440 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_70
timestamp 1623529830
transform 1 0 7544 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_82
timestamp 1623529830
transform 1 0 8648 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_94
timestamp 1623529830
transform 1 0 9752 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_106
timestamp 1623529830
transform 1 0 10856 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1623529830
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_115
timestamp 1623529830
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_127
timestamp 1623529830
transform 1 0 12788 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_139
timestamp 1623529830
transform 1 0 13892 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_151
timestamp 1623529830
transform 1 0 14996 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1623529830
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_163
timestamp 1623529830
transform 1 0 16100 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_172
timestamp 1623529830
transform 1 0 16928 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1623529830
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_196
timestamp 1623529830
transform 1 0 19136 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_Clk
timestamp 1623529830
transform -1 0 20240 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_204
timestamp 1623529830
transform 1 0 19872 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1623529830
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1623529830
transform 1 0 22080 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_220
timestamp 1623529830
transform 1 0 21344 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_229
timestamp 1623529830
transform 1 0 22172 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_241
timestamp 1623529830
transform 1 0 23276 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_253
timestamp 1623529830
transform 1 0 24380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_265
timestamp 1623529830
transform 1 0 25484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_277
timestamp 1623529830
transform 1 0 26588 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1623529830
transform 1 0 27324 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_286
timestamp 1623529830
transform 1 0 27416 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_298
timestamp 1623529830
transform 1 0 28520 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_310
timestamp 1623529830
transform 1 0 29624 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_322
timestamp 1623529830
transform 1 0 30728 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1623529830
transform 1 0 32568 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_334
timestamp 1623529830
transform 1 0 31832 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_343
timestamp 1623529830
transform 1 0 32660 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_355
timestamp 1623529830
transform 1 0 33764 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_367
timestamp 1623529830
transform 1 0 34868 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_379
timestamp 1623529830
transform 1 0 35972 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_391
timestamp 1623529830
transform 1 0 37076 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1623529830
transform -1 0 38824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1623529830
transform 1 0 37812 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_400
timestamp 1623529830
transform 1 0 37904 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_406
timestamp 1623529830
transform 1 0 38456 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1623529830
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1623529830
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1623529830
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1623529830
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1623529830
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_30
timestamp 1623529830
transform 1 0 3864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_42
timestamp 1623529830
transform 1 0 4968 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_54
timestamp 1623529830
transform 1 0 6072 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1623529830
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_66
timestamp 1623529830
transform 1 0 7176 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_78
timestamp 1623529830
transform 1 0 8280 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_87
timestamp 1623529830
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_99
timestamp 1623529830
transform 1 0 10212 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_111
timestamp 1623529830
transform 1 0 11316 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1623529830
transform 1 0 12420 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1623529830
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_135
timestamp 1623529830
transform 1 0 13524 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_144
timestamp 1623529830
transform 1 0 14352 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_156
timestamp 1623529830
transform 1 0 15456 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_168
timestamp 1623529830
transform 1 0 16560 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_180
timestamp 1623529830
transform 1 0 17664 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_192
timestamp 1623529830
transform 1 0 18768 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1623529830
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_201
timestamp 1623529830
transform 1 0 19596 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_213
timestamp 1623529830
transform 1 0 20700 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_225
timestamp 1623529830
transform 1 0 21804 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_237
timestamp 1623529830
transform 1 0 22908 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1623529830
transform 1 0 24748 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_249
timestamp 1623529830
transform 1 0 24012 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_258
timestamp 1623529830
transform 1 0 24840 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_270
timestamp 1623529830
transform 1 0 25944 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_282
timestamp 1623529830
transform 1 0 27048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_294
timestamp 1623529830
transform 1 0 28152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1623529830
transform 1 0 29992 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_306
timestamp 1623529830
transform 1 0 29256 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_315
timestamp 1623529830
transform 1 0 30084 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_327
timestamp 1623529830
transform 1 0 31188 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_339
timestamp 1623529830
transform 1 0 32292 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1623529830
transform 1 0 35236 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_351
timestamp 1623529830
transform 1 0 33396 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_363
timestamp 1623529830
transform 1 0 34500 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_372
timestamp 1623529830
transform 1 0 35328 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_384
timestamp 1623529830
transform 1 0 36432 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1623529830
transform -1 0 38824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_396
timestamp 1623529830
transform 1 0 37536 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_404
timestamp 1623529830
transform 1 0 38272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1623529830
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1623529830
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1623529830
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1623529830
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1623529830
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1623529830
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_51
timestamp 1623529830
transform 1 0 5796 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_58
timestamp 1623529830
transform 1 0 6440 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_70
timestamp 1623529830
transform 1 0 7544 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_82
timestamp 1623529830
transform 1 0 8648 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_94
timestamp 1623529830
transform 1 0 9752 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_106
timestamp 1623529830
transform 1 0 10856 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1623529830
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_115
timestamp 1623529830
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_127
timestamp 1623529830
transform 1 0 12788 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_139
timestamp 1623529830
transform 1 0 13892 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_151
timestamp 1623529830
transform 1 0 14996 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1623529830
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_163
timestamp 1623529830
transform 1 0 16100 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_172
timestamp 1623529830
transform 1 0 16928 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1623529830
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1623529830
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1623529830
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1623529830
transform 1 0 22080 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_220
timestamp 1623529830
transform 1 0 21344 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_229
timestamp 1623529830
transform 1 0 22172 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_241
timestamp 1623529830
transform 1 0 23276 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_253
timestamp 1623529830
transform 1 0 24380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_265
timestamp 1623529830
transform 1 0 25484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_277
timestamp 1623529830
transform 1 0 26588 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1623529830
transform 1 0 27324 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_286
timestamp 1623529830
transform 1 0 27416 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_298
timestamp 1623529830
transform 1 0 28520 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_310
timestamp 1623529830
transform 1 0 29624 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_322
timestamp 1623529830
transform 1 0 30728 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1623529830
transform 1 0 32568 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_334
timestamp 1623529830
transform 1 0 31832 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_343
timestamp 1623529830
transform 1 0 32660 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_355
timestamp 1623529830
transform 1 0 33764 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_367
timestamp 1623529830
transform 1 0 34868 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_379
timestamp 1623529830
transform 1 0 35972 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_391
timestamp 1623529830
transform 1 0 37076 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1623529830
transform -1 0 38824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1623529830
transform 1 0 37812 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_400
timestamp 1623529830
transform 1 0 37904 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_406
timestamp 1623529830
transform 1 0 38456 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1623529830
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1623529830
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1623529830
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1623529830
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1623529830
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1623529830
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1623529830
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1623529830
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_30
timestamp 1623529830
transform 1 0 3864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_42
timestamp 1623529830
transform 1 0 4968 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1623529830
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1623529830
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1623529830
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_54
timestamp 1623529830
transform 1 0 6072 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_51
timestamp 1623529830
transform 1 0 5796 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_58
timestamp 1623529830
transform 1 0 6440 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1623529830
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_66
timestamp 1623529830
transform 1 0 7176 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_78
timestamp 1623529830
transform 1 0 8280 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_87
timestamp 1623529830
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_70
timestamp 1623529830
transform 1 0 7544 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_82
timestamp 1623529830
transform 1 0 8648 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_99
timestamp 1623529830
transform 1 0 10212 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_94
timestamp 1623529830
transform 1 0 9752 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_106
timestamp 1623529830
transform 1 0 10856 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1623529830
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_111
timestamp 1623529830
transform 1 0 11316 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_123
timestamp 1623529830
transform 1 0 12420 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_115
timestamp 1623529830
transform 1 0 11684 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_127
timestamp 1623529830
transform 1 0 12788 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1623529830
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_135
timestamp 1623529830
transform 1 0 13524 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_144
timestamp 1623529830
transform 1 0 14352 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_139
timestamp 1623529830
transform 1 0 13892 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_151
timestamp 1623529830
transform 1 0 14996 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1623529830
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_156
timestamp 1623529830
transform 1 0 15456 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_168
timestamp 1623529830
transform 1 0 16560 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_163
timestamp 1623529830
transform 1 0 16100 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_172
timestamp 1623529830
transform 1 0 16928 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_180
timestamp 1623529830
transform 1 0 17664 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_192
timestamp 1623529830
transform 1 0 18768 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1623529830
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1623529830
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1623529830
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_201
timestamp 1623529830
transform 1 0 19596 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_213
timestamp 1623529830
transform 1 0 20700 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1623529830
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1623529830
transform 1 0 22080 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_225
timestamp 1623529830
transform 1 0 21804 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_237
timestamp 1623529830
transform 1 0 22908 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_220
timestamp 1623529830
transform 1 0 21344 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_229
timestamp 1623529830
transform 1 0 22172 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1623529830
transform 1 0 24748 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_249
timestamp 1623529830
transform 1 0 24012 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_258
timestamp 1623529830
transform 1 0 24840 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_241
timestamp 1623529830
transform 1 0 23276 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_253
timestamp 1623529830
transform 1 0 24380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_270
timestamp 1623529830
transform 1 0 25944 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_282
timestamp 1623529830
transform 1 0 27048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_265
timestamp 1623529830
transform 1 0 25484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_277
timestamp 1623529830
transform 1 0 26588 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1623529830
transform 1 0 27324 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_294
timestamp 1623529830
transform 1 0 28152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_286
timestamp 1623529830
transform 1 0 27416 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_298
timestamp 1623529830
transform 1 0 28520 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1623529830
transform 1 0 29992 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_306
timestamp 1623529830
transform 1 0 29256 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_315
timestamp 1623529830
transform 1 0 30084 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_327
timestamp 1623529830
transform 1 0 31188 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_310
timestamp 1623529830
transform 1 0 29624 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_322
timestamp 1623529830
transform 1 0 30728 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1623529830
transform 1 0 32568 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_339
timestamp 1623529830
transform 1 0 32292 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_334
timestamp 1623529830
transform 1 0 31832 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_343
timestamp 1623529830
transform 1 0 32660 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1623529830
transform 1 0 35236 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_351
timestamp 1623529830
transform 1 0 33396 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_363
timestamp 1623529830
transform 1 0 34500 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_355
timestamp 1623529830
transform 1 0 33764 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_367
timestamp 1623529830
transform 1 0 34868 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_372
timestamp 1623529830
transform 1 0 35328 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_384
timestamp 1623529830
transform 1 0 36432 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_379
timestamp 1623529830
transform 1 0 35972 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_391
timestamp 1623529830
transform 1 0 37076 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1623529830
transform -1 0 38824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1623529830
transform -1 0 38824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1623529830
transform 1 0 37812 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_396
timestamp 1623529830
transform 1 0 37536 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_404
timestamp 1623529830
transform 1 0 38272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_400
timestamp 1623529830
transform 1 0 37904 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_406
timestamp 1623529830
transform 1 0 38456 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1623529830
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1623529830
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1623529830
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1623529830
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1623529830
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_30
timestamp 1623529830
transform 1 0 3864 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_42
timestamp 1623529830
transform 1 0 4968 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_54
timestamp 1623529830
transform 1 0 6072 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1623529830
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_66
timestamp 1623529830
transform 1 0 7176 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_78
timestamp 1623529830
transform 1 0 8280 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_87
timestamp 1623529830
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_99
timestamp 1623529830
transform 1 0 10212 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_111
timestamp 1623529830
transform 1 0 11316 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_123
timestamp 1623529830
transform 1 0 12420 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1623529830
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_135
timestamp 1623529830
transform 1 0 13524 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_144
timestamp 1623529830
transform 1 0 14352 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_156
timestamp 1623529830
transform 1 0 15456 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_168
timestamp 1623529830
transform 1 0 16560 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_180
timestamp 1623529830
transform 1 0 17664 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_192
timestamp 1623529830
transform 1 0 18768 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfstp_1  _242_
timestamp 1623529830
transform 1 0 20884 0 -1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1623529830
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_201
timestamp 1623529830
transform 1 0 19596 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_213
timestamp 1623529830
transform 1 0 20700 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_236
timestamp 1623529830
transform 1 0 22816 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1623529830
transform 1 0 24748 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_248
timestamp 1623529830
transform 1 0 23920 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_256
timestamp 1623529830
transform 1 0 24656 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_258
timestamp 1623529830
transform 1 0 24840 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_270
timestamp 1623529830
transform 1 0 25944 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_282
timestamp 1623529830
transform 1 0 27048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_294
timestamp 1623529830
transform 1 0 28152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1623529830
transform 1 0 29992 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_306
timestamp 1623529830
transform 1 0 29256 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_315
timestamp 1623529830
transform 1 0 30084 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_327
timestamp 1623529830
transform 1 0 31188 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_339
timestamp 1623529830
transform 1 0 32292 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1623529830
transform 1 0 35236 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_351
timestamp 1623529830
transform 1 0 33396 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_363
timestamp 1623529830
transform 1 0 34500 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_372
timestamp 1623529830
transform 1 0 35328 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_384
timestamp 1623529830
transform 1 0 36432 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1623529830
transform -1 0 38824 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_396
timestamp 1623529830
transform 1 0 37536 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_404
timestamp 1623529830
transform 1 0 38272 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1623529830
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1623529830
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1623529830
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1623529830
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1623529830
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1623529830
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_51
timestamp 1623529830
transform 1 0 5796 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_58
timestamp 1623529830
transform 1 0 6440 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_70
timestamp 1623529830
transform 1 0 7544 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_82
timestamp 1623529830
transform 1 0 8648 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_94
timestamp 1623529830
transform 1 0 9752 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_106
timestamp 1623529830
transform 1 0 10856 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1623529830
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_115
timestamp 1623529830
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_127
timestamp 1623529830
transform 1 0 12788 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_139
timestamp 1623529830
transform 1 0 13892 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_151
timestamp 1623529830
transform 1 0 14996 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1623529830
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_163
timestamp 1623529830
transform 1 0 16100 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_172
timestamp 1623529830
transform 1 0 16928 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1623529830
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1623529830
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1623529830
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1623529830
transform 1 0 22080 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_220
timestamp 1623529830
transform 1 0 21344 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_229
timestamp 1623529830
transform 1 0 22172 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_241
timestamp 1623529830
transform 1 0 23276 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_253
timestamp 1623529830
transform 1 0 24380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_265
timestamp 1623529830
transform 1 0 25484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_277
timestamp 1623529830
transform 1 0 26588 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1623529830
transform 1 0 27324 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_286
timestamp 1623529830
transform 1 0 27416 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_298
timestamp 1623529830
transform 1 0 28520 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_310
timestamp 1623529830
transform 1 0 29624 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_322
timestamp 1623529830
transform 1 0 30728 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1623529830
transform 1 0 32568 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_334
timestamp 1623529830
transform 1 0 31832 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_343
timestamp 1623529830
transform 1 0 32660 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_355
timestamp 1623529830
transform 1 0 33764 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_367
timestamp 1623529830
transform 1 0 34868 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_379
timestamp 1623529830
transform 1 0 35972 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_391
timestamp 1623529830
transform 1 0 37076 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1623529830
transform -1 0 38824 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1623529830
transform 1 0 37812 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_400
timestamp 1623529830
transform 1 0 37904 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_406
timestamp 1623529830
transform 1 0 38456 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1623529830
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1623529830
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1623529830
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1623529830
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1623529830
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_30
timestamp 1623529830
transform 1 0 3864 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_42
timestamp 1623529830
transform 1 0 4968 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_54
timestamp 1623529830
transform 1 0 6072 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1623529830
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_66
timestamp 1623529830
transform 1 0 7176 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_78
timestamp 1623529830
transform 1 0 8280 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_87
timestamp 1623529830
transform 1 0 9108 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_99
timestamp 1623529830
transform 1 0 10212 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_111
timestamp 1623529830
transform 1 0 11316 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_123
timestamp 1623529830
transform 1 0 12420 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1623529830
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_135
timestamp 1623529830
transform 1 0 13524 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_144
timestamp 1623529830
transform 1 0 14352 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_156
timestamp 1623529830
transform 1 0 15456 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_168
timestamp 1623529830
transform 1 0 16560 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_180
timestamp 1623529830
transform 1 0 17664 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_192
timestamp 1623529830
transform 1 0 18768 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1623529830
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_201
timestamp 1623529830
transform 1 0 19596 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_213
timestamp 1623529830
transform 1 0 20700 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_225
timestamp 1623529830
transform 1 0 21804 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_237
timestamp 1623529830
transform 1 0 22908 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1623529830
transform 1 0 24748 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_249
timestamp 1623529830
transform 1 0 24012 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_258
timestamp 1623529830
transform 1 0 24840 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_270
timestamp 1623529830
transform 1 0 25944 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_282
timestamp 1623529830
transform 1 0 27048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_294
timestamp 1623529830
transform 1 0 28152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1623529830
transform 1 0 29992 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_306
timestamp 1623529830
transform 1 0 29256 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_315
timestamp 1623529830
transform 1 0 30084 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_327
timestamp 1623529830
transform 1 0 31188 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_339
timestamp 1623529830
transform 1 0 32292 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1623529830
transform 1 0 35236 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_351
timestamp 1623529830
transform 1 0 33396 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_363
timestamp 1623529830
transform 1 0 34500 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_372
timestamp 1623529830
transform 1 0 35328 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_384
timestamp 1623529830
transform 1 0 36432 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1623529830
transform -1 0 38824 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_396
timestamp 1623529830
transform 1 0 37536 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_404
timestamp 1623529830
transform 1 0 38272 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1623529830
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1623529830
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1623529830
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1623529830
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1623529830
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1623529830
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_51
timestamp 1623529830
transform 1 0 5796 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_58
timestamp 1623529830
transform 1 0 6440 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_70
timestamp 1623529830
transform 1 0 7544 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_82
timestamp 1623529830
transform 1 0 8648 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_94
timestamp 1623529830
transform 1 0 9752 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_106
timestamp 1623529830
transform 1 0 10856 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1623529830
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_115
timestamp 1623529830
transform 1 0 11684 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_127
timestamp 1623529830
transform 1 0 12788 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_139
timestamp 1623529830
transform 1 0 13892 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_151
timestamp 1623529830
transform 1 0 14996 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1623529830
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_163
timestamp 1623529830
transform 1 0 16100 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_172
timestamp 1623529830
transform 1 0 16928 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1623529830
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1623529830
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1623529830
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1623529830
transform 1 0 22080 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_220
timestamp 1623529830
transform 1 0 21344 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_229
timestamp 1623529830
transform 1 0 22172 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_241
timestamp 1623529830
transform 1 0 23276 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_253
timestamp 1623529830
transform 1 0 24380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_265
timestamp 1623529830
transform 1 0 25484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_277
timestamp 1623529830
transform 1 0 26588 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1623529830
transform 1 0 27324 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_286
timestamp 1623529830
transform 1 0 27416 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_298
timestamp 1623529830
transform 1 0 28520 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_310
timestamp 1623529830
transform 1 0 29624 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_322
timestamp 1623529830
transform 1 0 30728 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1623529830
transform 1 0 32568 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_334
timestamp 1623529830
transform 1 0 31832 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_343
timestamp 1623529830
transform 1 0 32660 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_355
timestamp 1623529830
transform 1 0 33764 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_367
timestamp 1623529830
transform 1 0 34868 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_379
timestamp 1623529830
transform 1 0 35972 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_391
timestamp 1623529830
transform 1 0 37076 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1623529830
transform -1 0 38824 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1623529830
transform 1 0 37812 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_400
timestamp 1623529830
transform 1 0 37904 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_406
timestamp 1623529830
transform 1 0 38456 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1623529830
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1623529830
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1623529830
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1623529830
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_27
timestamp 1623529830
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_30
timestamp 1623529830
transform 1 0 3864 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_42
timestamp 1623529830
transform 1 0 4968 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_54
timestamp 1623529830
transform 1 0 6072 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1623529830
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_66
timestamp 1623529830
transform 1 0 7176 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_78
timestamp 1623529830
transform 1 0 8280 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_87
timestamp 1623529830
transform 1 0 9108 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_99
timestamp 1623529830
transform 1 0 10212 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_111
timestamp 1623529830
transform 1 0 11316 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_123
timestamp 1623529830
transform 1 0 12420 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1623529830
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_135
timestamp 1623529830
transform 1 0 13524 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_144
timestamp 1623529830
transform 1 0 14352 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1623529830
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1623529830
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_180
timestamp 1623529830
transform 1 0 17664 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_192
timestamp 1623529830
transform 1 0 18768 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dfstp_1  _243_
timestamp 1623529830
transform -1 0 22080 0 -1 20128
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1623529830
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_201
timestamp 1623529830
transform 1 0 19596 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_228
timestamp 1623529830
transform 1 0 22080 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_240
timestamp 1623529830
transform 1 0 23184 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1623529830
transform 1 0 24748 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_252
timestamp 1623529830
transform 1 0 24288 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_256
timestamp 1623529830
transform 1 0 24656 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_258
timestamp 1623529830
transform 1 0 24840 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_270
timestamp 1623529830
transform 1 0 25944 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_282
timestamp 1623529830
transform 1 0 27048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_294
timestamp 1623529830
transform 1 0 28152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1623529830
transform 1 0 29992 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_306
timestamp 1623529830
transform 1 0 29256 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_315
timestamp 1623529830
transform 1 0 30084 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_327
timestamp 1623529830
transform 1 0 31188 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_339
timestamp 1623529830
transform 1 0 32292 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1623529830
transform 1 0 35236 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_351
timestamp 1623529830
transform 1 0 33396 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_363
timestamp 1623529830
transform 1 0 34500 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_372
timestamp 1623529830
transform 1 0 35328 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_384
timestamp 1623529830
transform 1 0 36432 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1623529830
transform -1 0 38824 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_396
timestamp 1623529830
transform 1 0 37536 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_404
timestamp 1623529830
transform 1 0 38272 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1623529830
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1623529830
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1623529830
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1623529830
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1623529830
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1623529830
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1623529830
transform 1 0 3772 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1623529830
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1623529830
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1623529830
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_30
timestamp 1623529830
transform 1 0 3864 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_42
timestamp 1623529830
transform 1 0 4968 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1623529830
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_51
timestamp 1623529830
transform 1 0 5796 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_58
timestamp 1623529830
transform 1 0 6440 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_54
timestamp 1623529830
transform 1 0 6072 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1623529830
transform 1 0 9016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_70
timestamp 1623529830
transform 1 0 7544 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_82
timestamp 1623529830
transform 1 0 8648 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_66
timestamp 1623529830
transform 1 0 7176 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_78
timestamp 1623529830
transform 1 0 8280 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_87
timestamp 1623529830
transform 1 0 9108 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_94
timestamp 1623529830
transform 1 0 9752 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_106
timestamp 1623529830
transform 1 0 10856 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_99
timestamp 1623529830
transform 1 0 10212 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1623529830
transform 1 0 11592 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_115
timestamp 1623529830
transform 1 0 11684 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_127
timestamp 1623529830
transform 1 0 12788 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_111
timestamp 1623529830
transform 1 0 11316 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_123
timestamp 1623529830
transform 1 0 12420 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1623529830
transform 1 0 14260 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_139
timestamp 1623529830
transform 1 0 13892 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_151
timestamp 1623529830
transform 1 0 14996 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_135
timestamp 1623529830
transform 1 0 13524 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_144
timestamp 1623529830
transform 1 0 14352 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1623529830
transform 1 0 16836 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_163
timestamp 1623529830
transform 1 0 16100 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_172
timestamp 1623529830
transform 1 0 16928 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_156
timestamp 1623529830
transform 1 0 15456 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_168
timestamp 1623529830
transform 1 0 16560 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _182_
timestamp 1623529830
transform 1 0 18860 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1623529830
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_196
timestamp 1623529830
transform 1 0 19136 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_180
timestamp 1623529830
transform 1 0 17664 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_192
timestamp 1623529830
transform 1 0 18768 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_196
timestamp 1623529830
transform 1 0 19136 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _244_
timestamp 1623529830
transform 1 0 19688 0 1 20128
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _245_
timestamp 1623529830
transform 1 0 19964 0 -1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1623529830
transform 1 0 19504 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_201
timestamp 1623529830
transform 1 0 19596 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1623529830
transform 1 0 22080 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_223
timestamp 1623529830
transform 1 0 21620 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_227
timestamp 1623529830
transform 1 0 21988 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_229
timestamp 1623529830
transform 1 0 22172 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_226
timestamp 1623529830
transform 1 0 21896 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_238
timestamp 1623529830
transform 1 0 23000 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1623529830
transform 1 0 24748 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_241
timestamp 1623529830
transform 1 0 23276 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_253
timestamp 1623529830
transform 1 0 24380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_250
timestamp 1623529830
transform 1 0 24104 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_256
timestamp 1623529830
transform 1 0 24656 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_258
timestamp 1623529830
transform 1 0 24840 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_265
timestamp 1623529830
transform 1 0 25484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_277
timestamp 1623529830
transform 1 0 26588 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_270
timestamp 1623529830
transform 1 0 25944 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_282
timestamp 1623529830
transform 1 0 27048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1623529830
transform 1 0 27324 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_286
timestamp 1623529830
transform 1 0 27416 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_298
timestamp 1623529830
transform 1 0 28520 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_294
timestamp 1623529830
transform 1 0 28152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1623529830
transform 1 0 29992 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_310
timestamp 1623529830
transform 1 0 29624 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_322
timestamp 1623529830
transform 1 0 30728 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_306
timestamp 1623529830
transform 1 0 29256 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_315
timestamp 1623529830
transform 1 0 30084 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_327
timestamp 1623529830
transform 1 0 31188 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1623529830
transform 1 0 32568 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_334
timestamp 1623529830
transform 1 0 31832 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_343
timestamp 1623529830
transform 1 0 32660 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_339
timestamp 1623529830
transform 1 0 32292 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1623529830
transform 1 0 35236 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_355
timestamp 1623529830
transform 1 0 33764 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_367
timestamp 1623529830
transform 1 0 34868 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_351
timestamp 1623529830
transform 1 0 33396 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_363
timestamp 1623529830
transform 1 0 34500 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_379
timestamp 1623529830
transform 1 0 35972 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_391
timestamp 1623529830
transform 1 0 37076 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_372
timestamp 1623529830
transform 1 0 35328 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_384
timestamp 1623529830
transform 1 0 36432 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1623529830
transform -1 0 38824 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1623529830
transform -1 0 38824 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1623529830
transform 1 0 37812 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_400
timestamp 1623529830
transform 1 0 37904 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_406
timestamp 1623529830
transform 1 0 38456 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_396
timestamp 1623529830
transform 1 0 37536 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_404
timestamp 1623529830
transform 1 0 38272 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1623529830
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1623529830
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1623529830
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1623529830
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1623529830
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1623529830
transform 1 0 6348 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_51
timestamp 1623529830
transform 1 0 5796 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_58
timestamp 1623529830
transform 1 0 6440 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_70
timestamp 1623529830
transform 1 0 7544 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_82
timestamp 1623529830
transform 1 0 8648 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1623529830
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_106
timestamp 1623529830
transform 1 0 10856 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1623529830
transform 1 0 11592 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_115
timestamp 1623529830
transform 1 0 11684 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_127
timestamp 1623529830
transform 1 0 12788 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_139
timestamp 1623529830
transform 1 0 13892 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_151
timestamp 1623529830
transform 1 0 14996 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1623529830
transform 1 0 16836 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_163
timestamp 1623529830
transform 1 0 16100 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_172
timestamp 1623529830
transform 1 0 16928 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfstp_1  _246_
timestamp 1623529830
transform 1 0 18676 0 1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_35_184
timestamp 1623529830
transform 1 0 18032 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_190
timestamp 1623529830
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_212
timestamp 1623529830
transform 1 0 20608 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1623529830
transform 1 0 22080 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_224
timestamp 1623529830
transform 1 0 21712 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_229
timestamp 1623529830
transform 1 0 22172 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_241
timestamp 1623529830
transform 1 0 23276 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_253
timestamp 1623529830
transform 1 0 24380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_265
timestamp 1623529830
transform 1 0 25484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_277
timestamp 1623529830
transform 1 0 26588 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1623529830
transform 1 0 27324 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_286
timestamp 1623529830
transform 1 0 27416 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_298
timestamp 1623529830
transform 1 0 28520 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_310
timestamp 1623529830
transform 1 0 29624 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_322
timestamp 1623529830
transform 1 0 30728 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1623529830
transform 1 0 32568 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_334
timestamp 1623529830
transform 1 0 31832 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_343
timestamp 1623529830
transform 1 0 32660 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_355
timestamp 1623529830
transform 1 0 33764 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_367
timestamp 1623529830
transform 1 0 34868 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_379
timestamp 1623529830
transform 1 0 35972 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_391
timestamp 1623529830
transform 1 0 37076 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1623529830
transform -1 0 38824 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1623529830
transform 1 0 37812 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_400
timestamp 1623529830
transform 1 0 37904 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_406
timestamp 1623529830
transform 1 0 38456 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1623529830
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1623529830
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1623529830
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1623529830
transform 1 0 3772 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1623529830
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_30
timestamp 1623529830
transform 1 0 3864 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_42
timestamp 1623529830
transform 1 0 4968 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_54
timestamp 1623529830
transform 1 0 6072 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1623529830
transform 1 0 9016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_66
timestamp 1623529830
transform 1 0 7176 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_78
timestamp 1623529830
transform 1 0 8280 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_87
timestamp 1623529830
transform 1 0 9108 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_99
timestamp 1623529830
transform 1 0 10212 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_111
timestamp 1623529830
transform 1 0 11316 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_123
timestamp 1623529830
transform 1 0 12420 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1623529830
transform 1 0 14260 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_135
timestamp 1623529830
transform 1 0 13524 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_144
timestamp 1623529830
transform 1 0 14352 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_156
timestamp 1623529830
transform 1 0 15456 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_168
timestamp 1623529830
transform 1 0 16560 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_180
timestamp 1623529830
transform 1 0 17664 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_192
timestamp 1623529830
transform 1 0 18768 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1623529830
transform 1 0 19504 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_201
timestamp 1623529830
transform 1 0 19596 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_213
timestamp 1623529830
transform 1 0 20700 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_225
timestamp 1623529830
transform 1 0 21804 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_237
timestamp 1623529830
transform 1 0 22908 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1623529830
transform 1 0 24748 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_249
timestamp 1623529830
transform 1 0 24012 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_258
timestamp 1623529830
transform 1 0 24840 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_270
timestamp 1623529830
transform 1 0 25944 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_282
timestamp 1623529830
transform 1 0 27048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_294
timestamp 1623529830
transform 1 0 28152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1623529830
transform 1 0 29992 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_306
timestamp 1623529830
transform 1 0 29256 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_315
timestamp 1623529830
transform 1 0 30084 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_327
timestamp 1623529830
transform 1 0 31188 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_339
timestamp 1623529830
transform 1 0 32292 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1623529830
transform 1 0 35236 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_351
timestamp 1623529830
transform 1 0 33396 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_363
timestamp 1623529830
transform 1 0 34500 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_372
timestamp 1623529830
transform 1 0 35328 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_384
timestamp 1623529830
transform 1 0 36432 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1623529830
transform -1 0 38824 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_396
timestamp 1623529830
transform 1 0 37536 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_404
timestamp 1623529830
transform 1 0 38272 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1623529830
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1623529830
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1623529830
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1623529830
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1623529830
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1623529830
transform 1 0 6348 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_51
timestamp 1623529830
transform 1 0 5796 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_58
timestamp 1623529830
transform 1 0 6440 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_70
timestamp 1623529830
transform 1 0 7544 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_82
timestamp 1623529830
transform 1 0 8648 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_94
timestamp 1623529830
transform 1 0 9752 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_106
timestamp 1623529830
transform 1 0 10856 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1623529830
transform 1 0 11592 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_115
timestamp 1623529830
transform 1 0 11684 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_127
timestamp 1623529830
transform 1 0 12788 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_139
timestamp 1623529830
transform 1 0 13892 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_151
timestamp 1623529830
transform 1 0 14996 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1623529830
transform 1 0 16836 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_163
timestamp 1623529830
transform 1 0 16100 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_172
timestamp 1623529830
transform 1 0 16928 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1623529830
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1623529830
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1623529830
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1623529830
transform 1 0 22080 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_220
timestamp 1623529830
transform 1 0 21344 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_229
timestamp 1623529830
transform 1 0 22172 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_241
timestamp 1623529830
transform 1 0 23276 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_253
timestamp 1623529830
transform 1 0 24380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_265
timestamp 1623529830
transform 1 0 25484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_277
timestamp 1623529830
transform 1 0 26588 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1623529830
transform 1 0 27324 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_286
timestamp 1623529830
transform 1 0 27416 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_298
timestamp 1623529830
transform 1 0 28520 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_310
timestamp 1623529830
transform 1 0 29624 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_322
timestamp 1623529830
transform 1 0 30728 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1623529830
transform 1 0 32568 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_334
timestamp 1623529830
transform 1 0 31832 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_343
timestamp 1623529830
transform 1 0 32660 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_355
timestamp 1623529830
transform 1 0 33764 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_367
timestamp 1623529830
transform 1 0 34868 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_379
timestamp 1623529830
transform 1 0 35972 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_391
timestamp 1623529830
transform 1 0 37076 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1623529830
transform -1 0 38824 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1623529830
transform 1 0 37812 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_400
timestamp 1623529830
transform 1 0 37904 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_406
timestamp 1623529830
transform 1 0 38456 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1623529830
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1623529830
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1623529830
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1623529830
transform 1 0 3772 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_27
timestamp 1623529830
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_30
timestamp 1623529830
transform 1 0 3864 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_42
timestamp 1623529830
transform 1 0 4968 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_54
timestamp 1623529830
transform 1 0 6072 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1623529830
transform 1 0 9016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_66
timestamp 1623529830
transform 1 0 7176 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_78
timestamp 1623529830
transform 1 0 8280 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_87
timestamp 1623529830
transform 1 0 9108 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_99
timestamp 1623529830
transform 1 0 10212 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_111
timestamp 1623529830
transform 1 0 11316 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_123
timestamp 1623529830
transform 1 0 12420 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1623529830
transform 1 0 14260 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_135
timestamp 1623529830
transform 1 0 13524 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_144
timestamp 1623529830
transform 1 0 14352 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_156
timestamp 1623529830
transform 1 0 15456 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_168
timestamp 1623529830
transform 1 0 16560 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_180
timestamp 1623529830
transform 1 0 17664 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_192
timestamp 1623529830
transform 1 0 18768 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1623529830
transform 1 0 19504 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_201
timestamp 1623529830
transform 1 0 19596 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_213
timestamp 1623529830
transform 1 0 20700 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_225
timestamp 1623529830
transform 1 0 21804 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_237
timestamp 1623529830
transform 1 0 22908 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1623529830
transform 1 0 24748 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_249
timestamp 1623529830
transform 1 0 24012 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_258
timestamp 1623529830
transform 1 0 24840 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_270
timestamp 1623529830
transform 1 0 25944 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_282
timestamp 1623529830
transform 1 0 27048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_294
timestamp 1623529830
transform 1 0 28152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1623529830
transform 1 0 29992 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_306
timestamp 1623529830
transform 1 0 29256 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_315
timestamp 1623529830
transform 1 0 30084 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_327
timestamp 1623529830
transform 1 0 31188 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_339
timestamp 1623529830
transform 1 0 32292 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1623529830
transform 1 0 35236 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_351
timestamp 1623529830
transform 1 0 33396 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_363
timestamp 1623529830
transform 1 0 34500 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_372
timestamp 1623529830
transform 1 0 35328 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_384
timestamp 1623529830
transform 1 0 36432 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1623529830
transform -1 0 38824 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_396
timestamp 1623529830
transform 1 0 37536 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_404
timestamp 1623529830
transform 1 0 38272 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1623529830
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1623529830
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1623529830
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1623529830
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1623529830
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1623529830
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1623529830
transform 1 0 3772 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1623529830
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1623529830
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_27
timestamp 1623529830
transform 1 0 3588 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_30
timestamp 1623529830
transform 1 0 3864 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_42
timestamp 1623529830
transform 1 0 4968 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1623529830
transform 1 0 6348 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_51
timestamp 1623529830
transform 1 0 5796 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_58
timestamp 1623529830
transform 1 0 6440 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_54
timestamp 1623529830
transform 1 0 6072 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1623529830
transform 1 0 9016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_70
timestamp 1623529830
transform 1 0 7544 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_82
timestamp 1623529830
transform 1 0 8648 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_66
timestamp 1623529830
transform 1 0 7176 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_78
timestamp 1623529830
transform 1 0 8280 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_87
timestamp 1623529830
transform 1 0 9108 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_94
timestamp 1623529830
transform 1 0 9752 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_106
timestamp 1623529830
transform 1 0 10856 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_99
timestamp 1623529830
transform 1 0 10212 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1623529830
transform 1 0 11592 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_115
timestamp 1623529830
transform 1 0 11684 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_127
timestamp 1623529830
transform 1 0 12788 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_111
timestamp 1623529830
transform 1 0 11316 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_123
timestamp 1623529830
transform 1 0 12420 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1623529830
transform 1 0 14260 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_139
timestamp 1623529830
transform 1 0 13892 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_151
timestamp 1623529830
transform 1 0 14996 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_135
timestamp 1623529830
transform 1 0 13524 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_144
timestamp 1623529830
transform 1 0 14352 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1623529830
transform 1 0 16836 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_163
timestamp 1623529830
transform 1 0 16100 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_172
timestamp 1623529830
transform 1 0 16928 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_156
timestamp 1623529830
transform 1 0 15456 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_168
timestamp 1623529830
transform 1 0 16560 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1623529830
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_196
timestamp 1623529830
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_180
timestamp 1623529830
transform 1 0 17664 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_192
timestamp 1623529830
transform 1 0 18768 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1623529830
transform 1 0 19504 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1623529830
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_201
timestamp 1623529830
transform 1 0 19596 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_213
timestamp 1623529830
transform 1 0 20700 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1623529830
transform 1 0 22080 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_220
timestamp 1623529830
transform 1 0 21344 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_229
timestamp 1623529830
transform 1 0 22172 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_225
timestamp 1623529830
transform 1 0 21804 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_237
timestamp 1623529830
transform 1 0 22908 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1623529830
transform 1 0 24748 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_241
timestamp 1623529830
transform 1 0 23276 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_253
timestamp 1623529830
transform 1 0 24380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_249
timestamp 1623529830
transform 1 0 24012 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_258
timestamp 1623529830
transform 1 0 24840 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_265
timestamp 1623529830
transform 1 0 25484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_277
timestamp 1623529830
transform 1 0 26588 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_270
timestamp 1623529830
transform 1 0 25944 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_282
timestamp 1623529830
transform 1 0 27048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1623529830
transform 1 0 27324 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_286
timestamp 1623529830
transform 1 0 27416 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_298
timestamp 1623529830
transform 1 0 28520 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_294
timestamp 1623529830
transform 1 0 28152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1623529830
transform 1 0 29992 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_310
timestamp 1623529830
transform 1 0 29624 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_322
timestamp 1623529830
transform 1 0 30728 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_306
timestamp 1623529830
transform 1 0 29256 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_315
timestamp 1623529830
transform 1 0 30084 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_327
timestamp 1623529830
transform 1 0 31188 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1623529830
transform 1 0 32568 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_334
timestamp 1623529830
transform 1 0 31832 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_343
timestamp 1623529830
transform 1 0 32660 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_339
timestamp 1623529830
transform 1 0 32292 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1623529830
transform 1 0 35236 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_355
timestamp 1623529830
transform 1 0 33764 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_367
timestamp 1623529830
transform 1 0 34868 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_351
timestamp 1623529830
transform 1 0 33396 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_363
timestamp 1623529830
transform 1 0 34500 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_379
timestamp 1623529830
transform 1 0 35972 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_391
timestamp 1623529830
transform 1 0 37076 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_372
timestamp 1623529830
transform 1 0 35328 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_384
timestamp 1623529830
transform 1 0 36432 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1623529830
transform -1 0 38824 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1623529830
transform -1 0 38824 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1623529830
transform 1 0 37812 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_400
timestamp 1623529830
transform 1 0 37904 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_406
timestamp 1623529830
transform 1 0 38456 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_396
timestamp 1623529830
transform 1 0 37536 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_404
timestamp 1623529830
transform 1 0 38272 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1623529830
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1623529830
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1623529830
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1623529830
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1623529830
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1623529830
transform 1 0 6348 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_51
timestamp 1623529830
transform 1 0 5796 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_58
timestamp 1623529830
transform 1 0 6440 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_70
timestamp 1623529830
transform 1 0 7544 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_82
timestamp 1623529830
transform 1 0 8648 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_94
timestamp 1623529830
transform 1 0 9752 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_106
timestamp 1623529830
transform 1 0 10856 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1623529830
transform 1 0 11592 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_115
timestamp 1623529830
transform 1 0 11684 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_127
timestamp 1623529830
transform 1 0 12788 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_139
timestamp 1623529830
transform 1 0 13892 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_151
timestamp 1623529830
transform 1 0 14996 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1623529830
transform 1 0 16836 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_163
timestamp 1623529830
transform 1 0 16100 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_172
timestamp 1623529830
transform 1 0 16928 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1623529830
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1623529830
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1623529830
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1623529830
transform 1 0 22080 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_220
timestamp 1623529830
transform 1 0 21344 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_229
timestamp 1623529830
transform 1 0 22172 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_241
timestamp 1623529830
transform 1 0 23276 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_253
timestamp 1623529830
transform 1 0 24380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_265
timestamp 1623529830
transform 1 0 25484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_277
timestamp 1623529830
transform 1 0 26588 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1623529830
transform 1 0 27324 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_286
timestamp 1623529830
transform 1 0 27416 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_298
timestamp 1623529830
transform 1 0 28520 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_310
timestamp 1623529830
transform 1 0 29624 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_322
timestamp 1623529830
transform 1 0 30728 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1623529830
transform 1 0 32568 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_334
timestamp 1623529830
transform 1 0 31832 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_343
timestamp 1623529830
transform 1 0 32660 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_355
timestamp 1623529830
transform 1 0 33764 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_367
timestamp 1623529830
transform 1 0 34868 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_379
timestamp 1623529830
transform 1 0 35972 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_391
timestamp 1623529830
transform 1 0 37076 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1623529830
transform -1 0 38824 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1623529830
transform 1 0 37812 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_400
timestamp 1623529830
transform 1 0 37904 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_406
timestamp 1623529830
transform 1 0 38456 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1623529830
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1623529830
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1623529830
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1623529830
transform 1 0 3772 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_27
timestamp 1623529830
transform 1 0 3588 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_30
timestamp 1623529830
transform 1 0 3864 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_42
timestamp 1623529830
transform 1 0 4968 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_54
timestamp 1623529830
transform 1 0 6072 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1623529830
transform 1 0 9016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_66
timestamp 1623529830
transform 1 0 7176 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_78
timestamp 1623529830
transform 1 0 8280 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_87
timestamp 1623529830
transform 1 0 9108 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_99
timestamp 1623529830
transform 1 0 10212 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_111
timestamp 1623529830
transform 1 0 11316 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_123
timestamp 1623529830
transform 1 0 12420 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1623529830
transform 1 0 14260 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_135
timestamp 1623529830
transform 1 0 13524 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_144
timestamp 1623529830
transform 1 0 14352 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1623529830
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1623529830
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_180
timestamp 1623529830
transform 1 0 17664 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_192
timestamp 1623529830
transform 1 0 18768 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1623529830
transform 1 0 19504 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_201
timestamp 1623529830
transform 1 0 19596 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_213
timestamp 1623529830
transform 1 0 20700 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_225
timestamp 1623529830
transform 1 0 21804 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_237
timestamp 1623529830
transform 1 0 22908 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1623529830
transform 1 0 24748 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_249
timestamp 1623529830
transform 1 0 24012 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_258
timestamp 1623529830
transform 1 0 24840 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_270
timestamp 1623529830
transform 1 0 25944 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_282
timestamp 1623529830
transform 1 0 27048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_294
timestamp 1623529830
transform 1 0 28152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1623529830
transform 1 0 29992 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_306
timestamp 1623529830
transform 1 0 29256 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_315
timestamp 1623529830
transform 1 0 30084 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_327
timestamp 1623529830
transform 1 0 31188 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_339
timestamp 1623529830
transform 1 0 32292 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1623529830
transform 1 0 35236 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_351
timestamp 1623529830
transform 1 0 33396 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_363
timestamp 1623529830
transform 1 0 34500 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_372
timestamp 1623529830
transform 1 0 35328 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_384
timestamp 1623529830
transform 1 0 36432 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1623529830
transform -1 0 38824 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_396
timestamp 1623529830
transform 1 0 37536 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_404
timestamp 1623529830
transform 1 0 38272 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1623529830
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1623529830
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1623529830
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1623529830
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1623529830
transform 1 0 4692 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1623529830
transform 1 0 6348 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_51
timestamp 1623529830
transform 1 0 5796 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_58
timestamp 1623529830
transform 1 0 6440 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_70
timestamp 1623529830
transform 1 0 7544 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_82
timestamp 1623529830
transform 1 0 8648 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_94
timestamp 1623529830
transform 1 0 9752 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_106
timestamp 1623529830
transform 1 0 10856 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1623529830
transform 1 0 11592 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_115
timestamp 1623529830
transform 1 0 11684 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_127
timestamp 1623529830
transform 1 0 12788 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_139
timestamp 1623529830
transform 1 0 13892 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_151
timestamp 1623529830
transform 1 0 14996 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1623529830
transform 1 0 16836 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_163
timestamp 1623529830
transform 1 0 16100 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_172
timestamp 1623529830
transform 1 0 16928 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_184
timestamp 1623529830
transform 1 0 18032 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_196
timestamp 1623529830
transform 1 0 19136 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_208
timestamp 1623529830
transform 1 0 20240 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1623529830
transform 1 0 22080 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_220
timestamp 1623529830
transform 1 0 21344 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_229
timestamp 1623529830
transform 1 0 22172 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_241
timestamp 1623529830
transform 1 0 23276 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_253
timestamp 1623529830
transform 1 0 24380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_265
timestamp 1623529830
transform 1 0 25484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_277
timestamp 1623529830
transform 1 0 26588 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1623529830
transform 1 0 27324 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_286
timestamp 1623529830
transform 1 0 27416 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_298
timestamp 1623529830
transform 1 0 28520 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_310
timestamp 1623529830
transform 1 0 29624 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_322
timestamp 1623529830
transform 1 0 30728 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1623529830
transform 1 0 32568 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_334
timestamp 1623529830
transform 1 0 31832 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_343
timestamp 1623529830
transform 1 0 32660 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_355
timestamp 1623529830
transform 1 0 33764 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_367
timestamp 1623529830
transform 1 0 34868 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_379
timestamp 1623529830
transform 1 0 35972 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_391
timestamp 1623529830
transform 1 0 37076 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1623529830
transform -1 0 38824 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1623529830
transform 1 0 37812 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_400
timestamp 1623529830
transform 1 0 37904 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_406
timestamp 1623529830
transform 1 0 38456 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1623529830
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1623529830
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1623529830
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1623529830
transform 1 0 3772 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_27
timestamp 1623529830
transform 1 0 3588 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_30
timestamp 1623529830
transform 1 0 3864 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_42
timestamp 1623529830
transform 1 0 4968 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_54
timestamp 1623529830
transform 1 0 6072 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1623529830
transform 1 0 9016 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_66
timestamp 1623529830
transform 1 0 7176 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_78
timestamp 1623529830
transform 1 0 8280 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_87
timestamp 1623529830
transform 1 0 9108 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_99
timestamp 1623529830
transform 1 0 10212 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_111
timestamp 1623529830
transform 1 0 11316 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_123
timestamp 1623529830
transform 1 0 12420 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1623529830
transform 1 0 14260 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_135
timestamp 1623529830
transform 1 0 13524 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_144
timestamp 1623529830
transform 1 0 14352 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_156
timestamp 1623529830
transform 1 0 15456 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_168
timestamp 1623529830
transform 1 0 16560 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_180
timestamp 1623529830
transform 1 0 17664 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_192
timestamp 1623529830
transform 1 0 18768 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1623529830
transform 1 0 19504 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_201
timestamp 1623529830
transform 1 0 19596 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_213
timestamp 1623529830
transform 1 0 20700 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_225
timestamp 1623529830
transform 1 0 21804 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_237
timestamp 1623529830
transform 1 0 22908 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1623529830
transform 1 0 24748 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_249
timestamp 1623529830
transform 1 0 24012 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_258
timestamp 1623529830
transform 1 0 24840 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_270
timestamp 1623529830
transform 1 0 25944 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_282
timestamp 1623529830
transform 1 0 27048 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_294
timestamp 1623529830
transform 1 0 28152 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1623529830
transform 1 0 29992 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_306
timestamp 1623529830
transform 1 0 29256 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_315
timestamp 1623529830
transform 1 0 30084 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_327
timestamp 1623529830
transform 1 0 31188 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_339
timestamp 1623529830
transform 1 0 32292 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1623529830
transform 1 0 35236 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_351
timestamp 1623529830
transform 1 0 33396 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_363
timestamp 1623529830
transform 1 0 34500 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_372
timestamp 1623529830
transform 1 0 35328 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_384
timestamp 1623529830
transform 1 0 36432 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1623529830
transform -1 0 38824 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_396
timestamp 1623529830
transform 1 0 37536 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_404
timestamp 1623529830
transform 1 0 38272 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1623529830
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1623529830
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1623529830
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1623529830
transform 1 0 3588 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1623529830
transform 1 0 4692 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1623529830
transform 1 0 6348 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_51
timestamp 1623529830
transform 1 0 5796 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_58
timestamp 1623529830
transform 1 0 6440 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_70
timestamp 1623529830
transform 1 0 7544 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_82
timestamp 1623529830
transform 1 0 8648 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_94
timestamp 1623529830
transform 1 0 9752 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_106
timestamp 1623529830
transform 1 0 10856 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1623529830
transform 1 0 11592 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_115
timestamp 1623529830
transform 1 0 11684 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_127
timestamp 1623529830
transform 1 0 12788 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_139
timestamp 1623529830
transform 1 0 13892 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_151
timestamp 1623529830
transform 1 0 14996 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1623529830
transform 1 0 16836 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_163
timestamp 1623529830
transform 1 0 16100 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_172
timestamp 1623529830
transform 1 0 16928 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_184
timestamp 1623529830
transform 1 0 18032 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_196
timestamp 1623529830
transform 1 0 19136 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_208
timestamp 1623529830
transform 1 0 20240 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1623529830
transform 1 0 22080 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_220
timestamp 1623529830
transform 1 0 21344 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_229
timestamp 1623529830
transform 1 0 22172 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_241
timestamp 1623529830
transform 1 0 23276 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_253
timestamp 1623529830
transform 1 0 24380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_265
timestamp 1623529830
transform 1 0 25484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_277
timestamp 1623529830
transform 1 0 26588 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1623529830
transform 1 0 27324 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_286
timestamp 1623529830
transform 1 0 27416 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_298
timestamp 1623529830
transform 1 0 28520 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_310
timestamp 1623529830
transform 1 0 29624 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_322
timestamp 1623529830
transform 1 0 30728 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1623529830
transform 1 0 32568 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_334
timestamp 1623529830
transform 1 0 31832 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_343
timestamp 1623529830
transform 1 0 32660 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_355
timestamp 1623529830
transform 1 0 33764 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_367
timestamp 1623529830
transform 1 0 34868 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_379
timestamp 1623529830
transform 1 0 35972 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_391
timestamp 1623529830
transform 1 0 37076 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1623529830
transform -1 0 38824 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1623529830
transform 1 0 37812 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_400
timestamp 1623529830
transform 1 0 37904 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_406
timestamp 1623529830
transform 1 0 38456 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1623529830
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1623529830
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1623529830
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1623529830
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1623529830
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1623529830
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1623529830
transform 1 0 3772 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_27
timestamp 1623529830
transform 1 0 3588 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_30
timestamp 1623529830
transform 1 0 3864 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_42
timestamp 1623529830
transform 1 0 4968 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1623529830
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1623529830
transform 1 0 4692 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1623529830
transform 1 0 6348 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_54
timestamp 1623529830
transform 1 0 6072 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_51
timestamp 1623529830
transform 1 0 5796 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_58
timestamp 1623529830
transform 1 0 6440 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1623529830
transform 1 0 9016 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_66
timestamp 1623529830
transform 1 0 7176 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_78
timestamp 1623529830
transform 1 0 8280 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_87
timestamp 1623529830
transform 1 0 9108 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_70
timestamp 1623529830
transform 1 0 7544 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_82
timestamp 1623529830
transform 1 0 8648 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_99
timestamp 1623529830
transform 1 0 10212 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_94
timestamp 1623529830
transform 1 0 9752 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_106
timestamp 1623529830
transform 1 0 10856 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1623529830
transform 1 0 11592 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_111
timestamp 1623529830
transform 1 0 11316 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_123
timestamp 1623529830
transform 1 0 12420 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_115
timestamp 1623529830
transform 1 0 11684 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_127
timestamp 1623529830
transform 1 0 12788 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1623529830
transform 1 0 14260 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_135
timestamp 1623529830
transform 1 0 13524 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_144
timestamp 1623529830
transform 1 0 14352 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_139
timestamp 1623529830
transform 1 0 13892 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_151
timestamp 1623529830
transform 1 0 14996 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1623529830
transform 1 0 16836 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_156
timestamp 1623529830
transform 1 0 15456 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_168
timestamp 1623529830
transform 1 0 16560 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_163
timestamp 1623529830
transform 1 0 16100 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_172
timestamp 1623529830
transform 1 0 16928 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_180
timestamp 1623529830
transform 1 0 17664 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_192
timestamp 1623529830
transform 1 0 18768 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_184
timestamp 1623529830
transform 1 0 18032 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_196
timestamp 1623529830
transform 1 0 19136 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1623529830
transform 1 0 19504 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_201
timestamp 1623529830
transform 1 0 19596 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_213
timestamp 1623529830
transform 1 0 20700 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_208
timestamp 1623529830
transform 1 0 20240 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1623529830
transform 1 0 22080 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_225
timestamp 1623529830
transform 1 0 21804 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_237
timestamp 1623529830
transform 1 0 22908 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_220
timestamp 1623529830
transform 1 0 21344 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_229
timestamp 1623529830
transform 1 0 22172 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1623529830
transform 1 0 24748 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_249
timestamp 1623529830
transform 1 0 24012 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_258
timestamp 1623529830
transform 1 0 24840 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_241
timestamp 1623529830
transform 1 0 23276 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_253
timestamp 1623529830
transform 1 0 24380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_270
timestamp 1623529830
transform 1 0 25944 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_282
timestamp 1623529830
transform 1 0 27048 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_265
timestamp 1623529830
transform 1 0 25484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_277
timestamp 1623529830
transform 1 0 26588 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1623529830
transform 1 0 27324 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_294
timestamp 1623529830
transform 1 0 28152 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_286
timestamp 1623529830
transform 1 0 27416 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_298
timestamp 1623529830
transform 1 0 28520 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1623529830
transform 1 0 29992 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_306
timestamp 1623529830
transform 1 0 29256 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_315
timestamp 1623529830
transform 1 0 30084 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_327
timestamp 1623529830
transform 1 0 31188 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_310
timestamp 1623529830
transform 1 0 29624 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_322
timestamp 1623529830
transform 1 0 30728 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1623529830
transform 1 0 32568 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_339
timestamp 1623529830
transform 1 0 32292 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_334
timestamp 1623529830
transform 1 0 31832 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_343
timestamp 1623529830
transform 1 0 32660 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1623529830
transform 1 0 35236 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_351
timestamp 1623529830
transform 1 0 33396 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_363
timestamp 1623529830
transform 1 0 34500 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_355
timestamp 1623529830
transform 1 0 33764 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_367
timestamp 1623529830
transform 1 0 34868 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_372
timestamp 1623529830
transform 1 0 35328 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_384
timestamp 1623529830
transform 1 0 36432 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_379
timestamp 1623529830
transform 1 0 35972 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_391
timestamp 1623529830
transform 1 0 37076 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1623529830
transform -1 0 38824 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1623529830
transform -1 0 38824 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1623529830
transform 1 0 37812 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_396
timestamp 1623529830
transform 1 0 37536 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_404
timestamp 1623529830
transform 1 0 38272 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_400
timestamp 1623529830
transform 1 0 37904 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_406
timestamp 1623529830
transform 1 0 38456 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1623529830
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1623529830
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1623529830
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1623529830
transform 1 0 3772 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_27
timestamp 1623529830
transform 1 0 3588 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_30
timestamp 1623529830
transform 1 0 3864 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_42
timestamp 1623529830
transform 1 0 4968 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_54
timestamp 1623529830
transform 1 0 6072 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1623529830
transform 1 0 9016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_66
timestamp 1623529830
transform 1 0 7176 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_78
timestamp 1623529830
transform 1 0 8280 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_87
timestamp 1623529830
transform 1 0 9108 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_99
timestamp 1623529830
transform 1 0 10212 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_111
timestamp 1623529830
transform 1 0 11316 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_123
timestamp 1623529830
transform 1 0 12420 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1623529830
transform 1 0 14260 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_135
timestamp 1623529830
transform 1 0 13524 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_144
timestamp 1623529830
transform 1 0 14352 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_156
timestamp 1623529830
transform 1 0 15456 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_168
timestamp 1623529830
transform 1 0 16560 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_180
timestamp 1623529830
transform 1 0 17664 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_192
timestamp 1623529830
transform 1 0 18768 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1623529830
transform 1 0 19504 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_201
timestamp 1623529830
transform 1 0 19596 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_213
timestamp 1623529830
transform 1 0 20700 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_225
timestamp 1623529830
transform 1 0 21804 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_237
timestamp 1623529830
transform 1 0 22908 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1623529830
transform 1 0 24748 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_249
timestamp 1623529830
transform 1 0 24012 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_258
timestamp 1623529830
transform 1 0 24840 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_270
timestamp 1623529830
transform 1 0 25944 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_282
timestamp 1623529830
transform 1 0 27048 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_294
timestamp 1623529830
transform 1 0 28152 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1623529830
transform 1 0 29992 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_306
timestamp 1623529830
transform 1 0 29256 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_315
timestamp 1623529830
transform 1 0 30084 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_327
timestamp 1623529830
transform 1 0 31188 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_339
timestamp 1623529830
transform 1 0 32292 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1623529830
transform 1 0 35236 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_351
timestamp 1623529830
transform 1 0 33396 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_363
timestamp 1623529830
transform 1 0 34500 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_372
timestamp 1623529830
transform 1 0 35328 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_384
timestamp 1623529830
transform 1 0 36432 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1623529830
transform -1 0 38824 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_396
timestamp 1623529830
transform 1 0 37536 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_404
timestamp 1623529830
transform 1 0 38272 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1623529830
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1623529830
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1623529830
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1623529830
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1623529830
transform 1 0 4692 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1623529830
transform 1 0 6348 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_51
timestamp 1623529830
transform 1 0 5796 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_58
timestamp 1623529830
transform 1 0 6440 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_70
timestamp 1623529830
transform 1 0 7544 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_82
timestamp 1623529830
transform 1 0 8648 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_94
timestamp 1623529830
transform 1 0 9752 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_106
timestamp 1623529830
transform 1 0 10856 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1623529830
transform 1 0 11592 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_115
timestamp 1623529830
transform 1 0 11684 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_127
timestamp 1623529830
transform 1 0 12788 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_139
timestamp 1623529830
transform 1 0 13892 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_151
timestamp 1623529830
transform 1 0 14996 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1623529830
transform 1 0 16836 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_163
timestamp 1623529830
transform 1 0 16100 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_172
timestamp 1623529830
transform 1 0 16928 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_184
timestamp 1623529830
transform 1 0 18032 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_196
timestamp 1623529830
transform 1 0 19136 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_208
timestamp 1623529830
transform 1 0 20240 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1623529830
transform 1 0 22080 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_220
timestamp 1623529830
transform 1 0 21344 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_229
timestamp 1623529830
transform 1 0 22172 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_241
timestamp 1623529830
transform 1 0 23276 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_253
timestamp 1623529830
transform 1 0 24380 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_265
timestamp 1623529830
transform 1 0 25484 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_277
timestamp 1623529830
transform 1 0 26588 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1623529830
transform 1 0 27324 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_286
timestamp 1623529830
transform 1 0 27416 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_298
timestamp 1623529830
transform 1 0 28520 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_310
timestamp 1623529830
transform 1 0 29624 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_322
timestamp 1623529830
transform 1 0 30728 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1623529830
transform 1 0 32568 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_334
timestamp 1623529830
transform 1 0 31832 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_343
timestamp 1623529830
transform 1 0 32660 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_355
timestamp 1623529830
transform 1 0 33764 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_367
timestamp 1623529830
transform 1 0 34868 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_379
timestamp 1623529830
transform 1 0 35972 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_391
timestamp 1623529830
transform 1 0 37076 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1623529830
transform -1 0 38824 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1623529830
transform 1 0 37812 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_400
timestamp 1623529830
transform 1 0 37904 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_406
timestamp 1623529830
transform 1 0 38456 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1623529830
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1623529830
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1623529830
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1623529830
transform 1 0 3772 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_27
timestamp 1623529830
transform 1 0 3588 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_30
timestamp 1623529830
transform 1 0 3864 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_42
timestamp 1623529830
transform 1 0 4968 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_54
timestamp 1623529830
transform 1 0 6072 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1623529830
transform 1 0 9016 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_66
timestamp 1623529830
transform 1 0 7176 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_78
timestamp 1623529830
transform 1 0 8280 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_87
timestamp 1623529830
transform 1 0 9108 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_99
timestamp 1623529830
transform 1 0 10212 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_111
timestamp 1623529830
transform 1 0 11316 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_123
timestamp 1623529830
transform 1 0 12420 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1623529830
transform 1 0 14260 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_135
timestamp 1623529830
transform 1 0 13524 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_144
timestamp 1623529830
transform 1 0 14352 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_156
timestamp 1623529830
transform 1 0 15456 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_168
timestamp 1623529830
transform 1 0 16560 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_180
timestamp 1623529830
transform 1 0 17664 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_192
timestamp 1623529830
transform 1 0 18768 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1623529830
transform 1 0 19504 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_201
timestamp 1623529830
transform 1 0 19596 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_213
timestamp 1623529830
transform 1 0 20700 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_225
timestamp 1623529830
transform 1 0 21804 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_237
timestamp 1623529830
transform 1 0 22908 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1623529830
transform 1 0 24748 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_249
timestamp 1623529830
transform 1 0 24012 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_258
timestamp 1623529830
transform 1 0 24840 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_270
timestamp 1623529830
transform 1 0 25944 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_282
timestamp 1623529830
transform 1 0 27048 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_294
timestamp 1623529830
transform 1 0 28152 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1623529830
transform 1 0 29992 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_306
timestamp 1623529830
transform 1 0 29256 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_315
timestamp 1623529830
transform 1 0 30084 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_327
timestamp 1623529830
transform 1 0 31188 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_339
timestamp 1623529830
transform 1 0 32292 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1623529830
transform 1 0 35236 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_351
timestamp 1623529830
transform 1 0 33396 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_363
timestamp 1623529830
transform 1 0 34500 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_372
timestamp 1623529830
transform 1 0 35328 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_384
timestamp 1623529830
transform 1 0 36432 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1623529830
transform -1 0 38824 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_396
timestamp 1623529830
transform 1 0 37536 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_404
timestamp 1623529830
transform 1 0 38272 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1623529830
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1623529830
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1623529830
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1623529830
transform 1 0 3588 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1623529830
transform 1 0 4692 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1623529830
transform 1 0 6348 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_51
timestamp 1623529830
transform 1 0 5796 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_58
timestamp 1623529830
transform 1 0 6440 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_70
timestamp 1623529830
transform 1 0 7544 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_82
timestamp 1623529830
transform 1 0 8648 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_94
timestamp 1623529830
transform 1 0 9752 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_106
timestamp 1623529830
transform 1 0 10856 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1623529830
transform 1 0 11592 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_115
timestamp 1623529830
transform 1 0 11684 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_127
timestamp 1623529830
transform 1 0 12788 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_139
timestamp 1623529830
transform 1 0 13892 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_151
timestamp 1623529830
transform 1 0 14996 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1623529830
transform 1 0 16836 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_163
timestamp 1623529830
transform 1 0 16100 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_172
timestamp 1623529830
transform 1 0 16928 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_184
timestamp 1623529830
transform 1 0 18032 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_196
timestamp 1623529830
transform 1 0 19136 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_208
timestamp 1623529830
transform 1 0 20240 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1623529830
transform 1 0 22080 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_220
timestamp 1623529830
transform 1 0 21344 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_229
timestamp 1623529830
transform 1 0 22172 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_241
timestamp 1623529830
transform 1 0 23276 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_253
timestamp 1623529830
transform 1 0 24380 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_265
timestamp 1623529830
transform 1 0 25484 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_277
timestamp 1623529830
transform 1 0 26588 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1623529830
transform 1 0 27324 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_286
timestamp 1623529830
transform 1 0 27416 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_298
timestamp 1623529830
transform 1 0 28520 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_310
timestamp 1623529830
transform 1 0 29624 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_322
timestamp 1623529830
transform 1 0 30728 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1623529830
transform 1 0 32568 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_334
timestamp 1623529830
transform 1 0 31832 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_343
timestamp 1623529830
transform 1 0 32660 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_355
timestamp 1623529830
transform 1 0 33764 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_367
timestamp 1623529830
transform 1 0 34868 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_379
timestamp 1623529830
transform 1 0 35972 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_391
timestamp 1623529830
transform 1 0 37076 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1623529830
transform -1 0 38824 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1623529830
transform 1 0 37812 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_400
timestamp 1623529830
transform 1 0 37904 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_406
timestamp 1623529830
transform 1 0 38456 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1623529830
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1623529830
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1623529830
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1623529830
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1623529830
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1623529830
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1623529830
transform 1 0 3772 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_27
timestamp 1623529830
transform 1 0 3588 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_30
timestamp 1623529830
transform 1 0 3864 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_42
timestamp 1623529830
transform 1 0 4968 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1623529830
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1623529830
transform 1 0 4692 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1623529830
transform 1 0 6348 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_54
timestamp 1623529830
transform 1 0 6072 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_51
timestamp 1623529830
transform 1 0 5796 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_58
timestamp 1623529830
transform 1 0 6440 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1623529830
transform 1 0 9016 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_66
timestamp 1623529830
transform 1 0 7176 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_78
timestamp 1623529830
transform 1 0 8280 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_87
timestamp 1623529830
transform 1 0 9108 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_70
timestamp 1623529830
transform 1 0 7544 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_82
timestamp 1623529830
transform 1 0 8648 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_99
timestamp 1623529830
transform 1 0 10212 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_94
timestamp 1623529830
transform 1 0 9752 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_106
timestamp 1623529830
transform 1 0 10856 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1623529830
transform 1 0 11592 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_111
timestamp 1623529830
transform 1 0 11316 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_123
timestamp 1623529830
transform 1 0 12420 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_115
timestamp 1623529830
transform 1 0 11684 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_127
timestamp 1623529830
transform 1 0 12788 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1623529830
transform 1 0 14260 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_135
timestamp 1623529830
transform 1 0 13524 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_144
timestamp 1623529830
transform 1 0 14352 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_139
timestamp 1623529830
transform 1 0 13892 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_151
timestamp 1623529830
transform 1 0 14996 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1623529830
transform 1 0 16836 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_156
timestamp 1623529830
transform 1 0 15456 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_168
timestamp 1623529830
transform 1 0 16560 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_163
timestamp 1623529830
transform 1 0 16100 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_172
timestamp 1623529830
transform 1 0 16928 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_180
timestamp 1623529830
transform 1 0 17664 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_192
timestamp 1623529830
transform 1 0 18768 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_184
timestamp 1623529830
transform 1 0 18032 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_196
timestamp 1623529830
transform 1 0 19136 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1623529830
transform 1 0 19504 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_201
timestamp 1623529830
transform 1 0 19596 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_213
timestamp 1623529830
transform 1 0 20700 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_208
timestamp 1623529830
transform 1 0 20240 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1623529830
transform 1 0 22080 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_225
timestamp 1623529830
transform 1 0 21804 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_237
timestamp 1623529830
transform 1 0 22908 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_220
timestamp 1623529830
transform 1 0 21344 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_229
timestamp 1623529830
transform 1 0 22172 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1623529830
transform 1 0 24748 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_249
timestamp 1623529830
transform 1 0 24012 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_258
timestamp 1623529830
transform 1 0 24840 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_241
timestamp 1623529830
transform 1 0 23276 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_253
timestamp 1623529830
transform 1 0 24380 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_270
timestamp 1623529830
transform 1 0 25944 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_282
timestamp 1623529830
transform 1 0 27048 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_265
timestamp 1623529830
transform 1 0 25484 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_277
timestamp 1623529830
transform 1 0 26588 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1623529830
transform 1 0 27324 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_294
timestamp 1623529830
transform 1 0 28152 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_286
timestamp 1623529830
transform 1 0 27416 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_298
timestamp 1623529830
transform 1 0 28520 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1623529830
transform 1 0 29992 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_306
timestamp 1623529830
transform 1 0 29256 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_315
timestamp 1623529830
transform 1 0 30084 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_327
timestamp 1623529830
transform 1 0 31188 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_310
timestamp 1623529830
transform 1 0 29624 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_322
timestamp 1623529830
transform 1 0 30728 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1623529830
transform 1 0 32568 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_339
timestamp 1623529830
transform 1 0 32292 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_334
timestamp 1623529830
transform 1 0 31832 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_343
timestamp 1623529830
transform 1 0 32660 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1623529830
transform 1 0 35236 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_351
timestamp 1623529830
transform 1 0 33396 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_363
timestamp 1623529830
transform 1 0 34500 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_355
timestamp 1623529830
transform 1 0 33764 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_367
timestamp 1623529830
transform 1 0 34868 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_372
timestamp 1623529830
transform 1 0 35328 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_384
timestamp 1623529830
transform 1 0 36432 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_379
timestamp 1623529830
transform 1 0 35972 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_391
timestamp 1623529830
transform 1 0 37076 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1623529830
transform -1 0 38824 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1623529830
transform -1 0 38824 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1623529830
transform 1 0 37812 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_396
timestamp 1623529830
transform 1 0 37536 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_404
timestamp 1623529830
transform 1 0 38272 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_400
timestamp 1623529830
transform 1 0 37904 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_406
timestamp 1623529830
transform 1 0 38456 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1623529830
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1623529830
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1623529830
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1623529830
transform 1 0 3772 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_27
timestamp 1623529830
transform 1 0 3588 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_30
timestamp 1623529830
transform 1 0 3864 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_42
timestamp 1623529830
transform 1 0 4968 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_54
timestamp 1623529830
transform 1 0 6072 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1623529830
transform 1 0 9016 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_66
timestamp 1623529830
transform 1 0 7176 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_78
timestamp 1623529830
transform 1 0 8280 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_87
timestamp 1623529830
transform 1 0 9108 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_99
timestamp 1623529830
transform 1 0 10212 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_111
timestamp 1623529830
transform 1 0 11316 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_123
timestamp 1623529830
transform 1 0 12420 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1623529830
transform 1 0 14260 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_135
timestamp 1623529830
transform 1 0 13524 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_144
timestamp 1623529830
transform 1 0 14352 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_156
timestamp 1623529830
transform 1 0 15456 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_168
timestamp 1623529830
transform 1 0 16560 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_180
timestamp 1623529830
transform 1 0 17664 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_192
timestamp 1623529830
transform 1 0 18768 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1623529830
transform 1 0 19504 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_201
timestamp 1623529830
transform 1 0 19596 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_213
timestamp 1623529830
transform 1 0 20700 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_225
timestamp 1623529830
transform 1 0 21804 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_237
timestamp 1623529830
transform 1 0 22908 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1623529830
transform 1 0 24748 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_249
timestamp 1623529830
transform 1 0 24012 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_258
timestamp 1623529830
transform 1 0 24840 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_270
timestamp 1623529830
transform 1 0 25944 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_282
timestamp 1623529830
transform 1 0 27048 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_294
timestamp 1623529830
transform 1 0 28152 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1623529830
transform 1 0 29992 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_306
timestamp 1623529830
transform 1 0 29256 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_315
timestamp 1623529830
transform 1 0 30084 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_327
timestamp 1623529830
transform 1 0 31188 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_339
timestamp 1623529830
transform 1 0 32292 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1623529830
transform 1 0 35236 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_351
timestamp 1623529830
transform 1 0 33396 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_363
timestamp 1623529830
transform 1 0 34500 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_372
timestamp 1623529830
transform 1 0 35328 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_384
timestamp 1623529830
transform 1 0 36432 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1623529830
transform -1 0 38824 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_396
timestamp 1623529830
transform 1 0 37536 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_404
timestamp 1623529830
transform 1 0 38272 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1623529830
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1623529830
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1623529830
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1623529830
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1623529830
transform 1 0 4692 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1623529830
transform 1 0 6348 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_51
timestamp 1623529830
transform 1 0 5796 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_58
timestamp 1623529830
transform 1 0 6440 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_70
timestamp 1623529830
transform 1 0 7544 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_82
timestamp 1623529830
transform 1 0 8648 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_94
timestamp 1623529830
transform 1 0 9752 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_106
timestamp 1623529830
transform 1 0 10856 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1623529830
transform 1 0 11592 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_115
timestamp 1623529830
transform 1 0 11684 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_127
timestamp 1623529830
transform 1 0 12788 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_139
timestamp 1623529830
transform 1 0 13892 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_151
timestamp 1623529830
transform 1 0 14996 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1623529830
transform 1 0 16836 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_163
timestamp 1623529830
transform 1 0 16100 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_172
timestamp 1623529830
transform 1 0 16928 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_184
timestamp 1623529830
transform 1 0 18032 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_196
timestamp 1623529830
transform 1 0 19136 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_208
timestamp 1623529830
transform 1 0 20240 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1623529830
transform 1 0 22080 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_220
timestamp 1623529830
transform 1 0 21344 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_229
timestamp 1623529830
transform 1 0 22172 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_241
timestamp 1623529830
transform 1 0 23276 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_253
timestamp 1623529830
transform 1 0 24380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_265
timestamp 1623529830
transform 1 0 25484 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_277
timestamp 1623529830
transform 1 0 26588 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1623529830
transform 1 0 27324 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_286
timestamp 1623529830
transform 1 0 27416 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_298
timestamp 1623529830
transform 1 0 28520 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_310
timestamp 1623529830
transform 1 0 29624 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_322
timestamp 1623529830
transform 1 0 30728 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1623529830
transform 1 0 32568 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_334
timestamp 1623529830
transform 1 0 31832 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_343
timestamp 1623529830
transform 1 0 32660 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_355
timestamp 1623529830
transform 1 0 33764 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_367
timestamp 1623529830
transform 1 0 34868 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_379
timestamp 1623529830
transform 1 0 35972 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_391
timestamp 1623529830
transform 1 0 37076 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1623529830
transform -1 0 38824 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1623529830
transform 1 0 37812 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_400
timestamp 1623529830
transform 1 0 37904 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_406
timestamp 1623529830
transform 1 0 38456 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1623529830
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1623529830
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1623529830
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1623529830
transform 1 0 3772 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_27
timestamp 1623529830
transform 1 0 3588 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_30
timestamp 1623529830
transform 1 0 3864 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_42
timestamp 1623529830
transform 1 0 4968 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_54
timestamp 1623529830
transform 1 0 6072 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1623529830
transform 1 0 9016 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_66
timestamp 1623529830
transform 1 0 7176 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_78
timestamp 1623529830
transform 1 0 8280 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_87
timestamp 1623529830
transform 1 0 9108 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_99
timestamp 1623529830
transform 1 0 10212 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_111
timestamp 1623529830
transform 1 0 11316 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_123
timestamp 1623529830
transform 1 0 12420 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1623529830
transform 1 0 14260 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_135
timestamp 1623529830
transform 1 0 13524 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_144
timestamp 1623529830
transform 1 0 14352 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_156
timestamp 1623529830
transform 1 0 15456 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_168
timestamp 1623529830
transform 1 0 16560 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_180
timestamp 1623529830
transform 1 0 17664 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_192
timestamp 1623529830
transform 1 0 18768 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1623529830
transform 1 0 19504 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_201
timestamp 1623529830
transform 1 0 19596 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_213
timestamp 1623529830
transform 1 0 20700 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_225
timestamp 1623529830
transform 1 0 21804 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_237
timestamp 1623529830
transform 1 0 22908 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1623529830
transform 1 0 24748 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_249
timestamp 1623529830
transform 1 0 24012 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_258
timestamp 1623529830
transform 1 0 24840 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_270
timestamp 1623529830
transform 1 0 25944 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_282
timestamp 1623529830
transform 1 0 27048 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_294
timestamp 1623529830
transform 1 0 28152 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1623529830
transform 1 0 29992 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_306
timestamp 1623529830
transform 1 0 29256 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_315
timestamp 1623529830
transform 1 0 30084 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_327
timestamp 1623529830
transform 1 0 31188 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_339
timestamp 1623529830
transform 1 0 32292 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1623529830
transform 1 0 35236 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_351
timestamp 1623529830
transform 1 0 33396 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_363
timestamp 1623529830
transform 1 0 34500 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_372
timestamp 1623529830
transform 1 0 35328 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_384
timestamp 1623529830
transform 1 0 36432 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1623529830
transform -1 0 38824 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_396
timestamp 1623529830
transform 1 0 37536 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_404
timestamp 1623529830
transform 1 0 38272 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1623529830
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1623529830
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1623529830
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1623529830
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1623529830
transform 1 0 4692 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1623529830
transform 1 0 6348 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_51
timestamp 1623529830
transform 1 0 5796 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_58
timestamp 1623529830
transform 1 0 6440 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_70
timestamp 1623529830
transform 1 0 7544 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_82
timestamp 1623529830
transform 1 0 8648 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_94
timestamp 1623529830
transform 1 0 9752 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_106
timestamp 1623529830
transform 1 0 10856 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1623529830
transform 1 0 11592 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_115
timestamp 1623529830
transform 1 0 11684 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_127
timestamp 1623529830
transform 1 0 12788 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_139
timestamp 1623529830
transform 1 0 13892 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_151
timestamp 1623529830
transform 1 0 14996 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1623529830
transform 1 0 16836 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_163
timestamp 1623529830
transform 1 0 16100 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_172
timestamp 1623529830
transform 1 0 16928 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_184
timestamp 1623529830
transform 1 0 18032 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_196
timestamp 1623529830
transform 1 0 19136 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_208
timestamp 1623529830
transform 1 0 20240 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1623529830
transform 1 0 22080 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_220
timestamp 1623529830
transform 1 0 21344 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_229
timestamp 1623529830
transform 1 0 22172 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_241
timestamp 1623529830
transform 1 0 23276 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_253
timestamp 1623529830
transform 1 0 24380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_265
timestamp 1623529830
transform 1 0 25484 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_277
timestamp 1623529830
transform 1 0 26588 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1623529830
transform 1 0 27324 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_286
timestamp 1623529830
transform 1 0 27416 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_298
timestamp 1623529830
transform 1 0 28520 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_310
timestamp 1623529830
transform 1 0 29624 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_322
timestamp 1623529830
transform 1 0 30728 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1623529830
transform 1 0 32568 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_334
timestamp 1623529830
transform 1 0 31832 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_343
timestamp 1623529830
transform 1 0 32660 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_355
timestamp 1623529830
transform 1 0 33764 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_367
timestamp 1623529830
transform 1 0 34868 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_379
timestamp 1623529830
transform 1 0 35972 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_391
timestamp 1623529830
transform 1 0 37076 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1623529830
transform -1 0 38824 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1623529830
transform 1 0 37812 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_400
timestamp 1623529830
transform 1 0 37904 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_406
timestamp 1623529830
transform 1 0 38456 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1623529830
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1623529830
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1623529830
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1623529830
transform 1 0 3772 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_27
timestamp 1623529830
transform 1 0 3588 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_30
timestamp 1623529830
transform 1 0 3864 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_42
timestamp 1623529830
transform 1 0 4968 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_54
timestamp 1623529830
transform 1 0 6072 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1623529830
transform 1 0 9016 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_66
timestamp 1623529830
transform 1 0 7176 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_78
timestamp 1623529830
transform 1 0 8280 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_87
timestamp 1623529830
transform 1 0 9108 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_99
timestamp 1623529830
transform 1 0 10212 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_111
timestamp 1623529830
transform 1 0 11316 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_123
timestamp 1623529830
transform 1 0 12420 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1623529830
transform 1 0 14260 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_135
timestamp 1623529830
transform 1 0 13524 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_144
timestamp 1623529830
transform 1 0 14352 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_156
timestamp 1623529830
transform 1 0 15456 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_168
timestamp 1623529830
transform 1 0 16560 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_180
timestamp 1623529830
transform 1 0 17664 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_192
timestamp 1623529830
transform 1 0 18768 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1623529830
transform 1 0 19504 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_201
timestamp 1623529830
transform 1 0 19596 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_213
timestamp 1623529830
transform 1 0 20700 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_225
timestamp 1623529830
transform 1 0 21804 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_237
timestamp 1623529830
transform 1 0 22908 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1623529830
transform 1 0 24748 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_249
timestamp 1623529830
transform 1 0 24012 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_258
timestamp 1623529830
transform 1 0 24840 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_270
timestamp 1623529830
transform 1 0 25944 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_282
timestamp 1623529830
transform 1 0 27048 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_294
timestamp 1623529830
transform 1 0 28152 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1623529830
transform 1 0 29992 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_306
timestamp 1623529830
transform 1 0 29256 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_315
timestamp 1623529830
transform 1 0 30084 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_327
timestamp 1623529830
transform 1 0 31188 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_339
timestamp 1623529830
transform 1 0 32292 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1623529830
transform 1 0 35236 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_351
timestamp 1623529830
transform 1 0 33396 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_363
timestamp 1623529830
transform 1 0 34500 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_372
timestamp 1623529830
transform 1 0 35328 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_384
timestamp 1623529830
transform 1 0 36432 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1623529830
transform -1 0 38824 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_396
timestamp 1623529830
transform 1 0 37536 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_404
timestamp 1623529830
transform 1 0 38272 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1623529830
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1623529830
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1623529830
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1623529830
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1623529830
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1623529830
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1623529830
transform 1 0 3772 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1623529830
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1623529830
transform 1 0 4692 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_27
timestamp 1623529830
transform 1 0 3588 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_30
timestamp 1623529830
transform 1 0 3864 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_42
timestamp 1623529830
transform 1 0 4968 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1623529830
transform 1 0 6348 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_51
timestamp 1623529830
transform 1 0 5796 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_58
timestamp 1623529830
transform 1 0 6440 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_54
timestamp 1623529830
transform 1 0 6072 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1623529830
transform 1 0 9016 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_70
timestamp 1623529830
transform 1 0 7544 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_82
timestamp 1623529830
transform 1 0 8648 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_66
timestamp 1623529830
transform 1 0 7176 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_78
timestamp 1623529830
transform 1 0 8280 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_87
timestamp 1623529830
transform 1 0 9108 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_94
timestamp 1623529830
transform 1 0 9752 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_106
timestamp 1623529830
transform 1 0 10856 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_99
timestamp 1623529830
transform 1 0 10212 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1623529830
transform 1 0 11592 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_115
timestamp 1623529830
transform 1 0 11684 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_127
timestamp 1623529830
transform 1 0 12788 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_111
timestamp 1623529830
transform 1 0 11316 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_123
timestamp 1623529830
transform 1 0 12420 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1623529830
transform 1 0 14260 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_139
timestamp 1623529830
transform 1 0 13892 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_151
timestamp 1623529830
transform 1 0 14996 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_135
timestamp 1623529830
transform 1 0 13524 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_144
timestamp 1623529830
transform 1 0 14352 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1623529830
transform 1 0 16836 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_163
timestamp 1623529830
transform 1 0 16100 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_172
timestamp 1623529830
transform 1 0 16928 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_156
timestamp 1623529830
transform 1 0 15456 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_168
timestamp 1623529830
transform 1 0 16560 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_184
timestamp 1623529830
transform 1 0 18032 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_196
timestamp 1623529830
transform 1 0 19136 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_180
timestamp 1623529830
transform 1 0 17664 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_192
timestamp 1623529830
transform 1 0 18768 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1623529830
transform 1 0 19504 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_208
timestamp 1623529830
transform 1 0 20240 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_201
timestamp 1623529830
transform 1 0 19596 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_213
timestamp 1623529830
transform 1 0 20700 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1623529830
transform 1 0 22080 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_220
timestamp 1623529830
transform 1 0 21344 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_229
timestamp 1623529830
transform 1 0 22172 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_225
timestamp 1623529830
transform 1 0 21804 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_237
timestamp 1623529830
transform 1 0 22908 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1623529830
transform 1 0 24748 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_241
timestamp 1623529830
transform 1 0 23276 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_253
timestamp 1623529830
transform 1 0 24380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_249
timestamp 1623529830
transform 1 0 24012 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_258
timestamp 1623529830
transform 1 0 24840 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_265
timestamp 1623529830
transform 1 0 25484 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_277
timestamp 1623529830
transform 1 0 26588 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_270
timestamp 1623529830
transform 1 0 25944 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_282
timestamp 1623529830
transform 1 0 27048 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1623529830
transform 1 0 27324 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_286
timestamp 1623529830
transform 1 0 27416 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_298
timestamp 1623529830
transform 1 0 28520 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_294
timestamp 1623529830
transform 1 0 28152 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1623529830
transform 1 0 29992 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_310
timestamp 1623529830
transform 1 0 29624 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_322
timestamp 1623529830
transform 1 0 30728 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_306
timestamp 1623529830
transform 1 0 29256 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_315
timestamp 1623529830
transform 1 0 30084 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_327
timestamp 1623529830
transform 1 0 31188 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1623529830
transform 1 0 32568 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_334
timestamp 1623529830
transform 1 0 31832 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_343
timestamp 1623529830
transform 1 0 32660 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_339
timestamp 1623529830
transform 1 0 32292 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1623529830
transform 1 0 35236 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_355
timestamp 1623529830
transform 1 0 33764 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_367
timestamp 1623529830
transform 1 0 34868 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_351
timestamp 1623529830
transform 1 0 33396 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_363
timestamp 1623529830
transform 1 0 34500 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_379
timestamp 1623529830
transform 1 0 35972 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_391
timestamp 1623529830
transform 1 0 37076 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_372
timestamp 1623529830
transform 1 0 35328 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_384
timestamp 1623529830
transform 1 0 36432 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1623529830
transform -1 0 38824 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1623529830
transform -1 0 38824 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1623529830
transform 1 0 37812 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_400
timestamp 1623529830
transform 1 0 37904 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_406
timestamp 1623529830
transform 1 0 38456 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_396
timestamp 1623529830
transform 1 0 37536 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_404
timestamp 1623529830
transform 1 0 38272 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1623529830
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1623529830
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1623529830
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1623529830
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1623529830
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1623529830
transform 1 0 6348 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_51
timestamp 1623529830
transform 1 0 5796 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_58
timestamp 1623529830
transform 1 0 6440 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_70
timestamp 1623529830
transform 1 0 7544 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_82
timestamp 1623529830
transform 1 0 8648 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_94
timestamp 1623529830
transform 1 0 9752 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_106
timestamp 1623529830
transform 1 0 10856 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1623529830
transform 1 0 11592 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_115
timestamp 1623529830
transform 1 0 11684 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_127
timestamp 1623529830
transform 1 0 12788 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_139
timestamp 1623529830
transform 1 0 13892 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_151
timestamp 1623529830
transform 1 0 14996 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1623529830
transform 1 0 16836 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_163
timestamp 1623529830
transform 1 0 16100 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_172
timestamp 1623529830
transform 1 0 16928 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_184
timestamp 1623529830
transform 1 0 18032 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_196
timestamp 1623529830
transform 1 0 19136 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_208
timestamp 1623529830
transform 1 0 20240 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1623529830
transform 1 0 22080 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_220
timestamp 1623529830
transform 1 0 21344 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_229
timestamp 1623529830
transform 1 0 22172 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_241
timestamp 1623529830
transform 1 0 23276 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_253
timestamp 1623529830
transform 1 0 24380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_265
timestamp 1623529830
transform 1 0 25484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_277
timestamp 1623529830
transform 1 0 26588 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1623529830
transform 1 0 27324 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_286
timestamp 1623529830
transform 1 0 27416 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_298
timestamp 1623529830
transform 1 0 28520 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_310
timestamp 1623529830
transform 1 0 29624 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_322
timestamp 1623529830
transform 1 0 30728 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1623529830
transform 1 0 32568 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_334
timestamp 1623529830
transform 1 0 31832 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_343
timestamp 1623529830
transform 1 0 32660 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_355
timestamp 1623529830
transform 1 0 33764 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_367
timestamp 1623529830
transform 1 0 34868 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_379
timestamp 1623529830
transform 1 0 35972 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_391
timestamp 1623529830
transform 1 0 37076 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1623529830
transform -1 0 38824 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1623529830
transform 1 0 37812 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_400
timestamp 1623529830
transform 1 0 37904 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_406
timestamp 1623529830
transform 1 0 38456 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1623529830
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1623529830
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1623529830
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1623529830
transform 1 0 3772 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_27
timestamp 1623529830
transform 1 0 3588 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_30
timestamp 1623529830
transform 1 0 3864 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_42
timestamp 1623529830
transform 1 0 4968 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_54
timestamp 1623529830
transform 1 0 6072 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1623529830
transform 1 0 9016 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_66
timestamp 1623529830
transform 1 0 7176 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_78
timestamp 1623529830
transform 1 0 8280 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_87
timestamp 1623529830
transform 1 0 9108 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_99
timestamp 1623529830
transform 1 0 10212 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_111
timestamp 1623529830
transform 1 0 11316 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_123
timestamp 1623529830
transform 1 0 12420 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1623529830
transform 1 0 14260 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_135
timestamp 1623529830
transform 1 0 13524 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_144
timestamp 1623529830
transform 1 0 14352 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_156
timestamp 1623529830
transform 1 0 15456 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_168
timestamp 1623529830
transform 1 0 16560 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_180
timestamp 1623529830
transform 1 0 17664 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_192
timestamp 1623529830
transform 1 0 18768 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1623529830
transform 1 0 19504 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_201
timestamp 1623529830
transform 1 0 19596 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_213
timestamp 1623529830
transform 1 0 20700 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_225
timestamp 1623529830
transform 1 0 21804 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_237
timestamp 1623529830
transform 1 0 22908 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1623529830
transform 1 0 24748 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_249
timestamp 1623529830
transform 1 0 24012 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_258
timestamp 1623529830
transform 1 0 24840 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_270
timestamp 1623529830
transform 1 0 25944 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_282
timestamp 1623529830
transform 1 0 27048 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_294
timestamp 1623529830
transform 1 0 28152 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1623529830
transform 1 0 29992 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_306
timestamp 1623529830
transform 1 0 29256 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_315
timestamp 1623529830
transform 1 0 30084 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_327
timestamp 1623529830
transform 1 0 31188 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_339
timestamp 1623529830
transform 1 0 32292 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1623529830
transform 1 0 35236 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_351
timestamp 1623529830
transform 1 0 33396 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_363
timestamp 1623529830
transform 1 0 34500 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_372
timestamp 1623529830
transform 1 0 35328 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_384
timestamp 1623529830
transform 1 0 36432 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1623529830
transform -1 0 38824 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_396
timestamp 1623529830
transform 1 0 37536 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_404
timestamp 1623529830
transform 1 0 38272 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1623529830
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1623529830
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1623529830
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1623529830
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1623529830
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1623529830
transform 1 0 6348 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_51
timestamp 1623529830
transform 1 0 5796 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_58
timestamp 1623529830
transform 1 0 6440 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_70
timestamp 1623529830
transform 1 0 7544 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_82
timestamp 1623529830
transform 1 0 8648 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_94
timestamp 1623529830
transform 1 0 9752 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_106
timestamp 1623529830
transform 1 0 10856 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1623529830
transform 1 0 11592 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_115
timestamp 1623529830
transform 1 0 11684 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_127
timestamp 1623529830
transform 1 0 12788 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_139
timestamp 1623529830
transform 1 0 13892 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_151
timestamp 1623529830
transform 1 0 14996 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1623529830
transform 1 0 16836 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_163
timestamp 1623529830
transform 1 0 16100 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_172
timestamp 1623529830
transform 1 0 16928 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_184
timestamp 1623529830
transform 1 0 18032 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_196
timestamp 1623529830
transform 1 0 19136 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 20240 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_212
timestamp 1623529830
transform 1 0 20608 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1623529830
transform 1 0 22080 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_224
timestamp 1623529830
transform 1 0 21712 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_229
timestamp 1623529830
transform 1 0 22172 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_241
timestamp 1623529830
transform 1 0 23276 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_253
timestamp 1623529830
transform 1 0 24380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_265
timestamp 1623529830
transform 1 0 25484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_277
timestamp 1623529830
transform 1 0 26588 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1623529830
transform 1 0 27324 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_286
timestamp 1623529830
transform 1 0 27416 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_298
timestamp 1623529830
transform 1 0 28520 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_310
timestamp 1623529830
transform 1 0 29624 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_322
timestamp 1623529830
transform 1 0 30728 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1623529830
transform 1 0 32568 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_334
timestamp 1623529830
transform 1 0 31832 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_343
timestamp 1623529830
transform 1 0 32660 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_355
timestamp 1623529830
transform 1 0 33764 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_367
timestamp 1623529830
transform 1 0 34868 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_379
timestamp 1623529830
transform 1 0 35972 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_391
timestamp 1623529830
transform 1 0 37076 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1623529830
transform -1 0 38824 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1623529830
transform 1 0 37812 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_400
timestamp 1623529830
transform 1 0 37904 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_406
timestamp 1623529830
transform 1 0 38456 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1623529830
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1623529830
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1623529830
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1623529830
transform 1 0 3772 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_27
timestamp 1623529830
transform 1 0 3588 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_30
timestamp 1623529830
transform 1 0 3864 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_42
timestamp 1623529830
transform 1 0 4968 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1623529830
transform 1 0 6440 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_54
timestamp 1623529830
transform 1 0 6072 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_59
timestamp 1623529830
transform 1 0 6532 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1623529830
transform 1 0 9108 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_71
timestamp 1623529830
transform 1 0 7636 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_83
timestamp 1623529830
transform 1 0 8740 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_88
timestamp 1623529830
transform 1 0 9200 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_100
timestamp 1623529830
transform 1 0 10304 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1623529830
transform 1 0 11776 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_112
timestamp 1623529830
transform 1 0 11408 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_117
timestamp 1623529830
transform 1 0 11868 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_129
timestamp 1623529830
transform 1 0 12972 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1623529830
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_141
timestamp 1623529830
transform 1 0 14076 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_146
timestamp 1623529830
transform 1 0 14536 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1623529830
transform 1 0 17112 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_158
timestamp 1623529830
transform 1 0 15640 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_170
timestamp 1623529830
transform 1 0 16744 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_175
timestamp 1623529830
transform 1 0 17204 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_187
timestamp 1623529830
transform 1 0 18308 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1623529830
transform 1 0 19780 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1623529830
transform 1 0 20424 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_199
timestamp 1623529830
transform 1 0 19412 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_204
timestamp 1623529830
transform 1 0 19872 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_218
timestamp 1623529830
transform 1 0 21160 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1623529830
transform 1 0 22448 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_230
timestamp 1623529830
transform 1 0 22264 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_233
timestamp 1623529830
transform 1 0 22540 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1623529830
transform 1 0 25116 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_245
timestamp 1623529830
transform 1 0 23644 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_257
timestamp 1623529830
transform 1 0 24748 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_262
timestamp 1623529830
transform 1 0 25208 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_274
timestamp 1623529830
transform 1 0 26312 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1623529830
transform 1 0 27784 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_286
timestamp 1623529830
transform 1 0 27416 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_291
timestamp 1623529830
transform 1 0 27876 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_303
timestamp 1623529830
transform 1 0 28980 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1623529830
transform 1 0 30452 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_315
timestamp 1623529830
transform 1 0 30084 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_320
timestamp 1623529830
transform 1 0 30544 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1623529830
transform 1 0 33120 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_332
timestamp 1623529830
transform 1 0 31648 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_344
timestamp 1623529830
transform 1 0 32752 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_349
timestamp 1623529830
transform 1 0 33212 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_361
timestamp 1623529830
transform 1 0 34316 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1623529830
transform 1 0 35788 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_373
timestamp 1623529830
transform 1 0 35420 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_378
timestamp 1623529830
transform 1 0 35880 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_390
timestamp 1623529830
transform 1 0 36984 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1623529830
transform -1 0 38824 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1623529830
transform 1 0 38456 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_402
timestamp 1623529830
transform 1 0 38088 0 -1 37536
box -38 -48 406 592
<< labels >>
rlabel metal2 s 19982 39200 20038 40000 6 ARstb
port 0 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 Clk
port 1 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 LFSR0out
port 2 nsew signal tristate
rlabel metal2 s 24398 0 24454 800 6 LFSR1in
port 3 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 LFSR1out
port 4 nsew signal tristate
rlabel metal2 s 37738 0 37794 800 6 io_oeb[0]
port 5 nsew signal tristate
rlabel metal2 s 28906 0 28962 800 6 io_oeb[1]
port 6 nsew signal tristate
rlabel metal2 s 19982 0 20038 800 6 io_oeb[2]
port 7 nsew signal tristate
rlabel metal2 s 11058 0 11114 800 6 io_oeb[3]
port 8 nsew signal tristate
rlabel metal2 s 2226 0 2282 800 6 io_oeb[4]
port 9 nsew signal tristate
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 10 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 11 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 12 nsew ground bidirectional
rlabel metal4 s 35588 2176 35908 37536 6 vccd2
port 13 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 37536 6 vccd2
port 14 nsew power bidirectional
rlabel metal4 s 20228 2176 20548 37536 6 vssd2
port 15 nsew ground bidirectional
rlabel metal4 s 36248 2176 36568 37536 6 vdda1
port 16 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 37536 6 vdda1
port 17 nsew power bidirectional
rlabel metal4 s 20888 2176 21208 37536 6 vssa1
port 18 nsew ground bidirectional
rlabel metal4 s 36908 2176 37228 37536 6 vdda2
port 19 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 37536 6 vdda2
port 20 nsew power bidirectional
rlabel metal4 s 21548 2176 21868 37536 6 vssa2
port 21 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
