magic
tech sky130A
magscale 1 2
timestamp 1624324453
<< nwell >>
rect 1066 36709 38862 37275
rect 1066 35621 38862 36187
rect 1066 34533 38862 35099
rect 1066 33445 38862 34011
rect 1066 32357 38862 32923
rect 1066 31269 38862 31835
rect 1066 30181 38862 30747
rect 1066 29093 38862 29659
rect 1066 28005 38862 28571
rect 1066 26917 38862 27483
rect 1066 25829 38862 26395
rect 1066 24741 38862 25307
rect 1066 23653 38862 24219
rect 1066 22565 38862 23131
rect 1066 21477 38862 22043
rect 1066 20389 38862 20955
rect 1066 19301 38862 19867
rect 1066 18213 38862 18779
rect 1066 17125 38862 17691
rect 1066 16037 38862 16603
rect 1066 14949 38862 15515
rect 1066 13861 38862 14427
rect 1066 12773 38862 13339
rect 1066 11685 38862 12251
rect 1066 10597 38862 11163
rect 1066 9509 38862 10075
rect 1066 8421 38862 8987
rect 1066 7333 38862 7899
rect 1066 6245 38862 6811
rect 1066 5157 38862 5723
rect 1066 4069 38862 4635
rect 1066 2981 38862 3547
rect 1066 2138 38862 2459
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 1104 960 38824 37584
<< metal2 >>
rect 19982 39200 20038 40000
rect 2226 0 2282 800
rect 6642 0 6698 800
rect 11058 0 11114 800
rect 15566 0 15622 800
rect 19982 0 20038 800
rect 24398 0 24454 800
rect 28906 0 28962 800
rect 33322 0 33378 800
rect 37738 0 37794 800
<< obsm2 >>
rect 2228 39144 19926 39200
rect 20094 39144 37792 39200
rect 2228 856 37792 39144
rect 2338 800 6586 856
rect 6754 800 11002 856
rect 11170 800 15510 856
rect 15678 800 19926 856
rect 20094 800 24342 856
rect 24510 800 28850 856
rect 29018 800 33266 856
rect 33434 800 37682 856
<< obsm3 >>
rect 4208 2143 35248 37569
<< metal4 >>
rect 4208 2128 4528 37584
rect 4868 2176 5188 37536
rect 5528 2176 5848 37536
rect 6188 2176 6508 37536
rect 19568 2128 19888 37584
rect 20228 2176 20548 37536
rect 20888 2176 21208 37536
rect 21548 2176 21868 37536
rect 34928 2128 35248 37584
rect 35588 2176 35908 37536
rect 36248 2176 36568 37536
rect 36908 2176 37228 37536
<< labels >>
rlabel metal2 s 19982 39200 20038 40000 6 ARstb
port 1 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 Clk
port 2 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 LFSR0out
port 3 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 LFSR1in
port 4 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 LFSR1out
port 5 nsew signal output
rlabel metal2 s 37738 0 37794 800 6 io_oeb[0]
port 6 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 io_oeb[1]
port 7 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 io_oeb[2]
port 8 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 io_oeb[3]
port 9 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 io_oeb[4]
port 10 nsew signal output
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 11 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 35588 2176 35908 37536 6 vccd2
port 14 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 37536 6 vccd2
port 15 nsew power bidirectional
rlabel metal4 s 20228 2176 20548 37536 6 vssd2
port 16 nsew ground bidirectional
rlabel metal4 s 36248 2176 36568 37536 6 vdda1
port 17 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 37536 6 vdda1
port 18 nsew power bidirectional
rlabel metal4 s 20888 2176 21208 37536 6 vssa1
port 19 nsew ground bidirectional
rlabel metal4 s 36908 2176 37228 37536 6 vdda2
port 20 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 37536 6 vdda2
port 21 nsew power bidirectional
rlabel metal4 s 21548 2176 21868 37536 6 vssa2
port 22 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 40000 40000
string LEFview TRUE
string GDS_FILE /project/openlane/lfsr32/runs/lfsr32/results/magic/lfsr32.gds
string GDS_END 785708
string GDS_START 107656
<< end >>

