magic
tech sky130A
magscale 1 2
timestamp 1624022286
<< locali >>
rect 25605 6647 25639 6749
<< viali >>
rect 38117 19873 38151 19907
rect 37933 19669 37967 19703
rect 33425 13277 33459 13311
rect 33793 13277 33827 13311
rect 31999 13141 32033 13175
rect 34851 12937 34885 12971
rect 30297 12801 30331 12835
rect 32091 12801 32125 12835
rect 33425 12801 33459 12835
rect 30665 12733 30699 12767
rect 33057 12733 33091 12767
rect 31217 12257 31251 12291
rect 32229 12257 32263 12291
rect 31861 12189 31895 12223
rect 33655 12053 33689 12087
rect 26801 11169 26835 11203
rect 33057 11169 33091 11203
rect 33425 11101 33459 11135
rect 26617 11033 26651 11067
rect 31631 11033 31665 11067
rect 26157 10693 26191 10727
rect 25513 10557 25547 10591
rect 26341 10557 26375 10591
rect 27997 10557 28031 10591
rect 25697 10421 25731 10455
rect 27813 10421 27847 10455
rect 31033 10217 31067 10251
rect 24133 10081 24167 10115
rect 25973 10081 26007 10115
rect 26617 10081 26651 10115
rect 27261 10081 27295 10115
rect 27721 10081 27755 10115
rect 28549 10081 28583 10115
rect 29009 10081 29043 10115
rect 30849 10081 30883 10115
rect 26433 9945 26467 9979
rect 28365 9945 28399 9979
rect 24317 9877 24351 9911
rect 25789 9877 25823 9911
rect 27077 9877 27111 9911
rect 27905 9877 27939 9911
rect 29193 9877 29227 9911
rect 24501 9605 24535 9639
rect 30389 9605 30423 9639
rect 24041 9469 24075 9503
rect 24685 9469 24719 9503
rect 27997 9469 28031 9503
rect 28641 9469 28675 9503
rect 29285 9469 29319 9503
rect 29937 9469 29971 9503
rect 30573 9469 30607 9503
rect 25145 9401 25179 9435
rect 23857 9333 23891 9367
rect 26433 9333 26467 9367
rect 27813 9333 27847 9367
rect 28457 9333 28491 9367
rect 29101 9333 29135 9367
rect 29745 9333 29779 9367
rect 22845 9129 22879 9163
rect 26709 9061 26743 9095
rect 23029 8993 23063 9027
rect 23673 8993 23707 9027
rect 24133 8993 24167 9027
rect 27445 8993 27479 9027
rect 28089 8993 28123 9027
rect 28917 8993 28951 9027
rect 29561 8993 29595 9027
rect 30665 8993 30699 9027
rect 31309 8993 31343 9027
rect 26985 8925 27019 8959
rect 28273 8857 28307 8891
rect 30481 8857 30515 8891
rect 31125 8857 31159 8891
rect 23489 8789 23523 8823
rect 24317 8789 24351 8823
rect 25237 8789 25271 8823
rect 27629 8789 27663 8823
rect 28733 8789 28767 8823
rect 29377 8789 29411 8823
rect 30205 8585 30239 8619
rect 31309 8585 31343 8619
rect 31861 8585 31895 8619
rect 24133 8517 24167 8551
rect 25145 8449 25179 8483
rect 26893 8449 26927 8483
rect 29285 8449 29319 8483
rect 22845 8381 22879 8415
rect 23673 8381 23707 8415
rect 24317 8381 24351 8415
rect 29561 8381 29595 8415
rect 30021 8381 30055 8415
rect 31401 8381 31435 8415
rect 32045 8381 32079 8415
rect 25421 8313 25455 8347
rect 23029 8245 23063 8279
rect 23489 8245 23523 8279
rect 27813 8245 27847 8279
rect 22569 8041 22603 8075
rect 28089 7973 28123 8007
rect 21289 7905 21323 7939
rect 22109 7905 22143 7939
rect 24317 7905 24351 7939
rect 30665 7905 30699 7939
rect 31301 7905 31335 7939
rect 31953 7905 31987 7939
rect 32597 7905 32631 7939
rect 33241 7905 33275 7939
rect 24041 7837 24075 7871
rect 25237 7837 25271 7871
rect 25513 7837 25547 7871
rect 27813 7837 27847 7871
rect 29561 7837 29595 7871
rect 21465 7769 21499 7803
rect 31769 7769 31803 7803
rect 33057 7769 33091 7803
rect 21925 7701 21959 7735
rect 26985 7701 27019 7735
rect 30481 7701 30515 7735
rect 31125 7701 31159 7735
rect 32413 7701 32447 7735
rect 20913 7497 20947 7531
rect 30665 7497 30699 7531
rect 31953 7497 31987 7531
rect 23581 7429 23615 7463
rect 23121 7361 23155 7395
rect 24593 7361 24627 7395
rect 20269 7293 20303 7327
rect 20845 7293 20879 7327
rect 21465 7293 21499 7327
rect 23305 7293 23339 7327
rect 23397 7293 23431 7327
rect 23673 7293 23707 7327
rect 29561 7293 29595 7327
rect 30021 7293 30055 7327
rect 30849 7293 30883 7327
rect 31493 7293 31527 7327
rect 32137 7293 32171 7327
rect 33241 7293 33275 7327
rect 33885 7293 33919 7327
rect 24869 7225 24903 7259
rect 29285 7225 29319 7259
rect 20085 7157 20119 7191
rect 21649 7157 21683 7191
rect 26341 7157 26375 7191
rect 27813 7157 27847 7191
rect 30205 7157 30239 7191
rect 31309 7157 31343 7191
rect 33057 7157 33091 7191
rect 33793 7157 33827 7191
rect 33517 6953 33551 6987
rect 25697 6817 25731 6851
rect 28641 6817 28675 6851
rect 29285 6817 29319 6851
rect 32689 6817 32723 6851
rect 33333 6817 33367 6851
rect 34161 6817 34195 6851
rect 34621 6817 34655 6851
rect 20361 6749 20395 6783
rect 20637 6749 20671 6783
rect 22569 6749 22603 6783
rect 22845 6749 22879 6783
rect 24317 6749 24351 6783
rect 25605 6749 25639 6783
rect 26341 6749 26375 6783
rect 27813 6749 27847 6783
rect 28089 6749 28123 6783
rect 32229 6749 32263 6783
rect 25881 6681 25915 6715
rect 29469 6681 29503 6715
rect 33977 6681 34011 6715
rect 22109 6613 22143 6647
rect 25605 6613 25639 6647
rect 28825 6613 28859 6647
rect 30481 6613 30515 6647
rect 31965 6613 31999 6647
rect 32873 6613 32907 6647
rect 34805 6613 34839 6647
rect 24685 6409 24719 6443
rect 34345 6409 34379 6443
rect 26893 6341 26927 6375
rect 30021 6341 30055 6375
rect 33701 6341 33735 6375
rect 22937 6273 22971 6307
rect 29561 6273 29595 6307
rect 31769 6273 31803 6307
rect 19441 6205 19475 6239
rect 19901 6205 19935 6239
rect 25145 6205 25179 6239
rect 27813 6205 27847 6239
rect 33241 6205 33275 6239
rect 33885 6205 33919 6239
rect 34537 6205 34571 6239
rect 34989 6205 35023 6239
rect 20177 6137 20211 6171
rect 23213 6137 23247 6171
rect 25421 6137 25455 6171
rect 28089 6137 28123 6171
rect 31493 6137 31527 6171
rect 19257 6069 19291 6103
rect 21649 6069 21683 6103
rect 33057 6069 33091 6103
rect 35081 6069 35115 6103
rect 18429 5865 18463 5899
rect 24317 5865 24351 5899
rect 30481 5865 30515 5899
rect 33977 5865 34011 5899
rect 35725 5865 35759 5899
rect 17601 5729 17635 5763
rect 18245 5729 18279 5763
rect 19073 5729 19107 5763
rect 22569 5729 22603 5763
rect 25513 5729 25547 5763
rect 25789 5729 25823 5763
rect 26525 5729 26559 5763
rect 29193 5729 29227 5763
rect 32873 5729 32907 5763
rect 33517 5729 33551 5763
rect 34161 5729 34195 5763
rect 34805 5729 34839 5763
rect 35909 5729 35943 5763
rect 20361 5661 20395 5695
rect 20637 5661 20671 5695
rect 22845 5661 22879 5695
rect 25421 5661 25455 5695
rect 25881 5661 25915 5695
rect 28457 5661 28491 5695
rect 28733 5661 28767 5695
rect 31953 5661 31987 5695
rect 32229 5661 32263 5695
rect 26341 5593 26375 5627
rect 34621 5593 34655 5627
rect 17417 5525 17451 5559
rect 18889 5525 18923 5559
rect 22109 5525 22143 5559
rect 25237 5525 25271 5559
rect 26985 5525 27019 5559
rect 29377 5525 29411 5559
rect 32689 5525 32723 5559
rect 33333 5525 33367 5559
rect 19177 5321 19211 5355
rect 21649 5321 21683 5355
rect 31769 5321 31803 5355
rect 35909 5321 35943 5355
rect 34805 5253 34839 5287
rect 36553 5253 36587 5287
rect 19441 5185 19475 5219
rect 19901 5185 19935 5219
rect 20177 5185 20211 5219
rect 24685 5185 24719 5219
rect 29285 5185 29319 5219
rect 29561 5185 29595 5219
rect 25145 5117 25179 5151
rect 30021 5117 30055 5151
rect 33057 5117 33091 5151
rect 35449 5117 35483 5151
rect 36093 5117 36127 5151
rect 36737 5117 36771 5151
rect 24409 5049 24443 5083
rect 25421 5049 25455 5083
rect 30297 5049 30331 5083
rect 33333 5049 33367 5083
rect 17693 4981 17727 5015
rect 22937 4981 22971 5015
rect 26893 4981 26927 5015
rect 27813 4981 27847 5015
rect 35265 4981 35299 5015
rect 35725 4777 35759 4811
rect 37657 4777 37691 4811
rect 25513 4709 25547 4743
rect 27721 4709 27755 4743
rect 30757 4709 30791 4743
rect 16681 4641 16715 4675
rect 17325 4641 17359 4675
rect 25237 4641 25271 4675
rect 30481 4641 30515 4675
rect 35909 4641 35943 4675
rect 36553 4641 36587 4675
rect 37197 4641 37231 4675
rect 37841 4641 37875 4675
rect 17601 4573 17635 4607
rect 20361 4573 20395 4607
rect 20637 4573 20671 4607
rect 22109 4573 22143 4607
rect 22569 4573 22603 4607
rect 22845 4573 22879 4607
rect 27445 4573 27479 4607
rect 29193 4573 29227 4607
rect 34161 4573 34195 4607
rect 34437 4573 34471 4607
rect 37013 4505 37047 4539
rect 16865 4437 16899 4471
rect 19073 4437 19107 4471
rect 24317 4437 24351 4471
rect 26985 4437 27019 4471
rect 32229 4437 32263 4471
rect 32689 4437 32723 4471
rect 36369 4437 36403 4471
rect 17956 4233 17990 4267
rect 20164 4233 20198 4267
rect 23200 4233 23234 4267
rect 25145 4233 25179 4267
rect 28070 4233 28104 4267
rect 29561 4233 29595 4267
rect 35265 4233 35299 4267
rect 19441 4097 19475 4131
rect 21649 4097 21683 4131
rect 22937 4097 22971 4131
rect 26617 4097 26651 4131
rect 26893 4097 26927 4131
rect 27813 4097 27847 4131
rect 30021 4097 30055 4131
rect 31493 4097 31527 4131
rect 15577 4029 15611 4063
rect 16221 4029 16255 4063
rect 17693 4029 17727 4063
rect 19901 4029 19935 4063
rect 31769 4029 31803 4063
rect 34805 4029 34839 4063
rect 35449 4029 35483 4063
rect 36093 4029 36127 4063
rect 36737 4029 36771 4063
rect 37381 4029 37415 4063
rect 34529 3961 34563 3995
rect 15761 3893 15795 3927
rect 16405 3893 16439 3927
rect 24685 3893 24719 3927
rect 33057 3893 33091 3927
rect 35909 3893 35943 3927
rect 36553 3893 36587 3927
rect 37197 3893 37231 3927
rect 19073 3689 19107 3723
rect 25237 3689 25271 3723
rect 28641 3689 28675 3723
rect 37473 3689 37507 3723
rect 37933 3689 37967 3723
rect 15393 3621 15427 3655
rect 20637 3621 20671 3655
rect 22845 3621 22879 3655
rect 25789 3621 25823 3655
rect 25881 3621 25915 3655
rect 27169 3621 27203 3655
rect 34161 3621 34195 3655
rect 36001 3621 36035 3655
rect 22569 3553 22603 3587
rect 25513 3553 25547 3587
rect 26893 3553 26927 3587
rect 29285 3553 29319 3587
rect 34437 3553 34471 3587
rect 35725 3553 35759 3587
rect 38117 3553 38151 3587
rect 15117 3485 15151 3519
rect 17325 3485 17359 3519
rect 17601 3485 17635 3519
rect 20361 3485 20395 3519
rect 24317 3485 24351 3519
rect 25421 3485 25455 3519
rect 31953 3485 31987 3519
rect 32229 3485 32263 3519
rect 16865 3417 16899 3451
rect 30481 3417 30515 3451
rect 22109 3349 22143 3383
rect 29101 3349 29135 3383
rect 32689 3349 32723 3383
rect 14105 3145 14139 3179
rect 17693 3145 17727 3179
rect 20164 3145 20198 3179
rect 21649 3145 21683 3179
rect 26893 3145 26927 3179
rect 33057 3145 33091 3179
rect 36921 3145 36955 3179
rect 16405 3077 16439 3111
rect 35265 3077 35299 3111
rect 22615 3009 22649 3043
rect 24041 3009 24075 3043
rect 24409 3009 24443 3043
rect 25145 3009 25179 3043
rect 25421 3009 25455 3043
rect 28641 3009 28675 3043
rect 29009 3009 29043 3043
rect 30941 3009 30975 3043
rect 31401 3009 31435 3043
rect 36461 3009 36495 3043
rect 14197 2941 14231 2975
rect 14657 2941 14691 2975
rect 19441 2941 19475 2975
rect 19901 2941 19935 2975
rect 27997 2941 28031 2975
rect 31309 2941 31343 2975
rect 34805 2941 34839 2975
rect 35449 2941 35483 2975
rect 35541 2941 35575 2975
rect 35817 2941 35851 2975
rect 36369 2941 36403 2975
rect 36645 2941 36679 2975
rect 36737 2941 36771 2975
rect 14933 2873 14967 2907
rect 19165 2873 19199 2907
rect 31033 2873 31067 2907
rect 34529 2873 34563 2907
rect 35909 2873 35943 2907
rect 28181 2805 28215 2839
rect 30435 2805 30469 2839
rect 31585 2805 31619 2839
rect 16037 2601 16071 2635
rect 16497 2601 16531 2635
rect 19349 2601 19383 2635
rect 22017 2601 22051 2635
rect 24685 2601 24719 2635
rect 30021 2601 30055 2635
rect 30941 2601 30975 2635
rect 35357 2601 35391 2635
rect 15117 2533 15151 2567
rect 17877 2533 17911 2567
rect 23213 2533 23247 2567
rect 27077 2533 27111 2567
rect 32413 2533 32447 2567
rect 33885 2533 33919 2567
rect 36461 2533 36495 2567
rect 13185 2465 13219 2499
rect 13829 2465 13863 2499
rect 15853 2465 15887 2499
rect 16681 2465 16715 2499
rect 20269 2465 20303 2499
rect 22937 2465 22971 2499
rect 27353 2465 27387 2499
rect 28273 2465 28307 2499
rect 32689 2465 32723 2499
rect 33609 2465 33643 2499
rect 37197 2465 37231 2499
rect 37841 2465 37875 2499
rect 17601 2397 17635 2431
rect 20545 2397 20579 2431
rect 25605 2397 25639 2431
rect 28549 2397 28583 2431
rect 14933 2329 14967 2363
rect 36277 2329 36311 2363
rect 37657 2329 37691 2363
rect 13369 2261 13403 2295
rect 14013 2261 14047 2295
rect 37013 2261 37047 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 38824 37562
rect 1104 37488 38824 37510
rect 1104 37018 38824 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 38824 37018
rect 1104 36944 38824 36966
rect 1104 36474 38824 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 38824 36474
rect 1104 36400 38824 36422
rect 1104 35930 38824 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 38824 35930
rect 1104 35856 38824 35878
rect 1104 35386 38824 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 38824 35386
rect 1104 35312 38824 35334
rect 1104 34842 38824 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 38824 34842
rect 1104 34768 38824 34790
rect 1104 34298 38824 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 38824 34298
rect 1104 34224 38824 34246
rect 1104 33754 38824 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 38824 33754
rect 1104 33680 38824 33702
rect 1104 33210 38824 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 38824 33210
rect 1104 33136 38824 33158
rect 1104 32666 38824 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 38824 32666
rect 1104 32592 38824 32614
rect 1104 32122 38824 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 38824 32122
rect 1104 32048 38824 32070
rect 1104 31578 38824 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 38824 31578
rect 1104 31504 38824 31526
rect 1104 31034 38824 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 38824 31034
rect 1104 30960 38824 30982
rect 1104 30490 38824 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 38824 30490
rect 1104 30416 38824 30438
rect 1104 29946 38824 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 38824 29946
rect 1104 29872 38824 29894
rect 1104 29402 38824 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 38824 29402
rect 1104 29328 38824 29350
rect 1104 28858 38824 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 38824 28858
rect 1104 28784 38824 28806
rect 1104 28314 38824 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 38824 28314
rect 1104 28240 38824 28262
rect 1104 27770 38824 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 38824 27770
rect 1104 27696 38824 27718
rect 1104 27226 38824 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 38824 27226
rect 1104 27152 38824 27174
rect 1104 26682 38824 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 38824 26682
rect 1104 26608 38824 26630
rect 1104 26138 38824 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 38824 26138
rect 1104 26064 38824 26086
rect 1104 25594 38824 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 38824 25594
rect 1104 25520 38824 25542
rect 1104 25050 38824 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 38824 25050
rect 1104 24976 38824 24998
rect 1104 24506 38824 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 38824 24506
rect 1104 24432 38824 24454
rect 1104 23962 38824 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 38824 23962
rect 1104 23888 38824 23910
rect 1104 23418 38824 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 38824 23418
rect 1104 23344 38824 23366
rect 1104 22874 38824 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 38824 22874
rect 1104 22800 38824 22822
rect 1104 22330 38824 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 38824 22330
rect 1104 22256 38824 22278
rect 1104 21786 38824 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 38824 21786
rect 1104 21712 38824 21734
rect 1104 21242 38824 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 38824 21242
rect 1104 21168 38824 21190
rect 1104 20698 38824 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 38824 20698
rect 1104 20624 38824 20646
rect 1104 20154 38824 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 38824 20154
rect 1104 20080 38824 20102
rect 38102 19904 38108 19916
rect 38063 19876 38108 19904
rect 38102 19864 38108 19876
rect 38160 19864 38166 19916
rect 35250 19660 35256 19712
rect 35308 19700 35314 19712
rect 37921 19703 37979 19709
rect 37921 19700 37933 19703
rect 35308 19672 37933 19700
rect 35308 19660 35314 19672
rect 37921 19669 37933 19672
rect 37967 19669 37979 19703
rect 37921 19663 37979 19669
rect 1104 19610 38824 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 38824 19610
rect 1104 19536 38824 19558
rect 1104 19066 38824 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 38824 19066
rect 1104 18992 38824 19014
rect 1104 18522 38824 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 38824 18522
rect 1104 18448 38824 18470
rect 1104 17978 38824 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 38824 17978
rect 1104 17904 38824 17926
rect 1104 17434 38824 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 38824 17434
rect 1104 17360 38824 17382
rect 1104 16890 38824 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 38824 16890
rect 1104 16816 38824 16838
rect 1104 16346 38824 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 38824 16346
rect 1104 16272 38824 16294
rect 1104 15802 38824 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 38824 15802
rect 1104 15728 38824 15750
rect 1104 15258 38824 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 38824 15258
rect 1104 15184 38824 15206
rect 1104 14714 38824 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 38824 14714
rect 1104 14640 38824 14662
rect 1104 14170 38824 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 38824 14170
rect 1104 14096 38824 14118
rect 1104 13626 38824 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 38824 13626
rect 1104 13552 38824 13574
rect 35250 13512 35256 13524
rect 33060 13484 35256 13512
rect 33060 13456 33088 13484
rect 35250 13472 35256 13484
rect 35308 13472 35314 13524
rect 33042 13404 33048 13456
rect 33100 13404 33106 13456
rect 33410 13308 33416 13320
rect 33371 13280 33416 13308
rect 33410 13268 33416 13280
rect 33468 13268 33474 13320
rect 33781 13311 33839 13317
rect 33781 13277 33793 13311
rect 33827 13277 33839 13311
rect 33781 13271 33839 13277
rect 31987 13175 32045 13181
rect 31987 13141 31999 13175
rect 32033 13172 32045 13175
rect 32214 13172 32220 13184
rect 32033 13144 32220 13172
rect 32033 13141 32045 13144
rect 31987 13135 32045 13141
rect 32214 13132 32220 13144
rect 32272 13132 32278 13184
rect 32950 13132 32956 13184
rect 33008 13172 33014 13184
rect 33796 13172 33824 13271
rect 33008 13144 33824 13172
rect 33008 13132 33014 13144
rect 1104 13082 38824 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 38824 13082
rect 1104 13008 38824 13030
rect 33410 12928 33416 12980
rect 33468 12968 33474 12980
rect 34839 12971 34897 12977
rect 34839 12968 34851 12971
rect 33468 12940 34851 12968
rect 33468 12928 33474 12940
rect 34839 12937 34851 12940
rect 34885 12937 34897 12971
rect 34839 12931 34897 12937
rect 30285 12835 30343 12841
rect 30285 12801 30297 12835
rect 30331 12832 30343 12835
rect 31846 12832 31852 12844
rect 30331 12804 31852 12832
rect 30331 12801 30343 12804
rect 30285 12795 30343 12801
rect 31846 12792 31852 12804
rect 31904 12792 31910 12844
rect 32079 12835 32137 12841
rect 32079 12801 32091 12835
rect 32125 12832 32137 12835
rect 33413 12835 33471 12841
rect 33413 12832 33425 12835
rect 32125 12804 33425 12832
rect 32125 12801 32137 12804
rect 32079 12795 32137 12801
rect 33413 12801 33425 12804
rect 33459 12801 33471 12835
rect 33413 12795 33471 12801
rect 30650 12764 30656 12776
rect 30611 12736 30656 12764
rect 30650 12724 30656 12736
rect 30708 12724 30714 12776
rect 31864 12764 31892 12792
rect 32950 12764 32956 12776
rect 31864 12736 32956 12764
rect 32950 12724 32956 12736
rect 33008 12764 33014 12776
rect 33045 12767 33103 12773
rect 33045 12764 33057 12767
rect 33008 12736 33057 12764
rect 33008 12724 33014 12736
rect 33045 12733 33057 12736
rect 33091 12733 33103 12767
rect 33045 12727 33103 12733
rect 35250 12696 35256 12708
rect 31680 12628 31708 12682
rect 34454 12668 35256 12696
rect 35250 12656 35256 12668
rect 35308 12656 35314 12708
rect 32674 12628 32680 12640
rect 31680 12600 32680 12628
rect 32674 12588 32680 12600
rect 32732 12628 32738 12640
rect 33042 12628 33048 12640
rect 32732 12600 33048 12628
rect 32732 12588 32738 12600
rect 33042 12588 33048 12600
rect 33100 12588 33106 12640
rect 1104 12538 38824 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 38824 12538
rect 1104 12464 38824 12486
rect 33042 12316 33048 12368
rect 33100 12316 33106 12368
rect 30650 12248 30656 12300
rect 30708 12288 30714 12300
rect 31205 12291 31263 12297
rect 31205 12288 31217 12291
rect 30708 12260 31217 12288
rect 30708 12248 30714 12260
rect 31205 12257 31217 12260
rect 31251 12257 31263 12291
rect 32214 12288 32220 12300
rect 32175 12260 32220 12288
rect 31205 12251 31263 12257
rect 32214 12248 32220 12260
rect 32272 12248 32278 12300
rect 31846 12220 31852 12232
rect 31807 12192 31852 12220
rect 31846 12180 31852 12192
rect 31904 12180 31910 12232
rect 33042 12044 33048 12096
rect 33100 12084 33106 12096
rect 33643 12087 33701 12093
rect 33643 12084 33655 12087
rect 33100 12056 33655 12084
rect 33100 12044 33106 12056
rect 33643 12053 33655 12056
rect 33689 12053 33701 12087
rect 33643 12047 33701 12053
rect 1104 11994 38824 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 38824 11994
rect 1104 11920 38824 11942
rect 1104 11450 38824 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 38824 11450
rect 1104 11376 38824 11398
rect 32674 11228 32680 11280
rect 32732 11228 32738 11280
rect 26789 11203 26847 11209
rect 26789 11169 26801 11203
rect 26835 11200 26847 11203
rect 27706 11200 27712 11212
rect 26835 11172 27712 11200
rect 26835 11169 26847 11172
rect 26789 11163 26847 11169
rect 27706 11160 27712 11172
rect 27764 11160 27770 11212
rect 33042 11200 33048 11212
rect 33003 11172 33048 11200
rect 33042 11160 33048 11172
rect 33100 11160 33106 11212
rect 31846 11092 31852 11144
rect 31904 11132 31910 11144
rect 33413 11135 33471 11141
rect 33413 11132 33425 11135
rect 31904 11104 33425 11132
rect 31904 11092 31910 11104
rect 33413 11101 33425 11104
rect 33459 11101 33471 11135
rect 33413 11095 33471 11101
rect 23658 11024 23664 11076
rect 23716 11064 23722 11076
rect 26605 11067 26663 11073
rect 26605 11064 26617 11067
rect 23716 11036 26617 11064
rect 23716 11024 23722 11036
rect 26605 11033 26617 11036
rect 26651 11033 26663 11067
rect 26605 11027 26663 11033
rect 31386 11024 31392 11076
rect 31444 11064 31450 11076
rect 31619 11067 31677 11073
rect 31619 11064 31631 11067
rect 31444 11036 31631 11064
rect 31444 11024 31450 11036
rect 31619 11033 31631 11036
rect 31665 11033 31677 11067
rect 31619 11027 31677 11033
rect 1104 10906 38824 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 38824 10906
rect 1104 10832 38824 10854
rect 24118 10684 24124 10736
rect 24176 10724 24182 10736
rect 26145 10727 26203 10733
rect 26145 10724 26157 10727
rect 24176 10696 26157 10724
rect 24176 10684 24182 10696
rect 26145 10693 26157 10696
rect 26191 10693 26203 10727
rect 26145 10687 26203 10693
rect 27246 10656 27252 10668
rect 25516 10628 27252 10656
rect 25516 10597 25544 10628
rect 27246 10616 27252 10628
rect 27304 10616 27310 10668
rect 25501 10591 25559 10597
rect 25501 10557 25513 10591
rect 25547 10557 25559 10591
rect 25501 10551 25559 10557
rect 26329 10591 26387 10597
rect 26329 10557 26341 10591
rect 26375 10588 26387 10591
rect 27890 10588 27896 10600
rect 26375 10560 27896 10588
rect 26375 10557 26387 10560
rect 26329 10551 26387 10557
rect 27890 10548 27896 10560
rect 27948 10548 27954 10600
rect 27985 10591 28043 10597
rect 27985 10557 27997 10591
rect 28031 10588 28043 10591
rect 30834 10588 30840 10600
rect 28031 10560 30840 10588
rect 28031 10557 28043 10560
rect 27985 10551 28043 10557
rect 30834 10548 30840 10560
rect 30892 10548 30898 10600
rect 31018 10520 31024 10532
rect 25700 10492 31024 10520
rect 25700 10461 25728 10492
rect 31018 10480 31024 10492
rect 31076 10480 31082 10532
rect 25685 10455 25743 10461
rect 25685 10421 25697 10455
rect 25731 10421 25743 10455
rect 27798 10452 27804 10464
rect 27759 10424 27804 10452
rect 25685 10415 25743 10421
rect 27798 10412 27804 10424
rect 27856 10412 27862 10464
rect 1104 10362 38824 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 38824 10362
rect 1104 10288 38824 10310
rect 31021 10251 31079 10257
rect 31021 10217 31033 10251
rect 31067 10248 31079 10251
rect 31846 10248 31852 10260
rect 31067 10220 31852 10248
rect 31067 10217 31079 10220
rect 31021 10211 31079 10217
rect 31846 10208 31852 10220
rect 31904 10208 31910 10260
rect 28902 10180 28908 10192
rect 27264 10152 28908 10180
rect 22830 10072 22836 10124
rect 22888 10112 22894 10124
rect 24121 10115 24179 10121
rect 24121 10112 24133 10115
rect 22888 10084 24133 10112
rect 22888 10072 22894 10084
rect 24121 10081 24133 10084
rect 24167 10081 24179 10115
rect 24121 10075 24179 10081
rect 25866 10072 25872 10124
rect 25924 10112 25930 10124
rect 27264 10121 27292 10152
rect 28902 10140 28908 10152
rect 28960 10140 28966 10192
rect 25961 10115 26019 10121
rect 25961 10112 25973 10115
rect 25924 10084 25973 10112
rect 25924 10072 25930 10084
rect 25961 10081 25973 10084
rect 26007 10081 26019 10115
rect 25961 10075 26019 10081
rect 26605 10115 26663 10121
rect 26605 10081 26617 10115
rect 26651 10081 26663 10115
rect 26605 10075 26663 10081
rect 27249 10115 27307 10121
rect 27249 10081 27261 10115
rect 27295 10081 27307 10115
rect 27706 10112 27712 10124
rect 27667 10084 27712 10112
rect 27249 10075 27307 10081
rect 26620 10044 26648 10075
rect 27706 10072 27712 10084
rect 27764 10072 27770 10124
rect 28537 10115 28595 10121
rect 28537 10081 28549 10115
rect 28583 10081 28595 10115
rect 28537 10075 28595 10081
rect 28997 10115 29055 10121
rect 28997 10081 29009 10115
rect 29043 10112 29055 10115
rect 30834 10112 30840 10124
rect 29043 10084 30052 10112
rect 30795 10084 30840 10112
rect 29043 10081 29055 10084
rect 28997 10075 29055 10081
rect 28074 10044 28080 10056
rect 26620 10016 28080 10044
rect 28074 10004 28080 10016
rect 28132 10004 28138 10056
rect 28552 10044 28580 10075
rect 29914 10044 29920 10056
rect 28552 10016 29920 10044
rect 29914 10004 29920 10016
rect 29972 10004 29978 10056
rect 30024 10044 30052 10084
rect 30834 10072 30840 10084
rect 30892 10072 30898 10124
rect 31202 10044 31208 10056
rect 30024 10016 31208 10044
rect 31202 10004 31208 10016
rect 31260 10004 31266 10056
rect 24946 9936 24952 9988
rect 25004 9976 25010 9988
rect 26421 9979 26479 9985
rect 26421 9976 26433 9979
rect 25004 9948 26433 9976
rect 25004 9936 25010 9948
rect 26421 9945 26433 9948
rect 26467 9945 26479 9979
rect 26421 9939 26479 9945
rect 26694 9936 26700 9988
rect 26752 9976 26758 9988
rect 28353 9979 28411 9985
rect 28353 9976 28365 9979
rect 26752 9948 28365 9976
rect 26752 9936 26758 9948
rect 28353 9945 28365 9948
rect 28399 9945 28411 9979
rect 28353 9939 28411 9945
rect 24302 9908 24308 9920
rect 24263 9880 24308 9908
rect 24302 9868 24308 9880
rect 24360 9868 24366 9920
rect 25774 9908 25780 9920
rect 25735 9880 25780 9908
rect 25774 9868 25780 9880
rect 25832 9868 25838 9920
rect 26326 9868 26332 9920
rect 26384 9908 26390 9920
rect 27065 9911 27123 9917
rect 27065 9908 27077 9911
rect 26384 9880 27077 9908
rect 26384 9868 26390 9880
rect 27065 9877 27077 9880
rect 27111 9877 27123 9911
rect 27065 9871 27123 9877
rect 27893 9911 27951 9917
rect 27893 9877 27905 9911
rect 27939 9908 27951 9911
rect 29086 9908 29092 9920
rect 27939 9880 29092 9908
rect 27939 9877 27951 9880
rect 27893 9871 27951 9877
rect 29086 9868 29092 9880
rect 29144 9868 29150 9920
rect 29181 9911 29239 9917
rect 29181 9877 29193 9911
rect 29227 9908 29239 9911
rect 30650 9908 30656 9920
rect 29227 9880 30656 9908
rect 29227 9877 29239 9880
rect 29181 9871 29239 9877
rect 30650 9868 30656 9880
rect 30708 9868 30714 9920
rect 1104 9818 38824 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 38824 9818
rect 1104 9744 38824 9766
rect 16114 9664 16120 9716
rect 16172 9704 16178 9716
rect 25774 9704 25780 9716
rect 16172 9676 25780 9704
rect 16172 9664 16178 9676
rect 25774 9664 25780 9676
rect 25832 9664 25838 9716
rect 23106 9596 23112 9648
rect 23164 9636 23170 9648
rect 24489 9639 24547 9645
rect 24489 9636 24501 9639
rect 23164 9608 24501 9636
rect 23164 9596 23170 9608
rect 24489 9605 24501 9608
rect 24535 9605 24547 9639
rect 24489 9599 24547 9605
rect 28718 9596 28724 9648
rect 28776 9636 28782 9648
rect 30377 9639 30435 9645
rect 30377 9636 30389 9639
rect 28776 9608 30389 9636
rect 28776 9596 28782 9608
rect 30377 9605 30389 9608
rect 30423 9605 30435 9639
rect 30377 9599 30435 9605
rect 27522 9528 27528 9580
rect 27580 9568 27586 9580
rect 32030 9568 32036 9580
rect 27580 9540 29408 9568
rect 27580 9528 27586 9540
rect 22922 9460 22928 9512
rect 22980 9500 22986 9512
rect 24029 9503 24087 9509
rect 24029 9500 24041 9503
rect 22980 9472 24041 9500
rect 22980 9460 22986 9472
rect 24029 9469 24041 9472
rect 24075 9469 24087 9503
rect 24670 9500 24676 9512
rect 24631 9472 24676 9500
rect 24029 9463 24087 9469
rect 24670 9460 24676 9472
rect 24728 9500 24734 9512
rect 25866 9500 25872 9512
rect 24728 9472 25872 9500
rect 24728 9460 24734 9472
rect 25866 9460 25872 9472
rect 25924 9460 25930 9512
rect 27614 9460 27620 9512
rect 27672 9500 27678 9512
rect 27985 9503 28043 9509
rect 27985 9500 27997 9503
rect 27672 9472 27997 9500
rect 27672 9460 27678 9472
rect 27985 9469 27997 9472
rect 28031 9469 28043 9503
rect 27985 9463 28043 9469
rect 28629 9503 28687 9509
rect 28629 9469 28641 9503
rect 28675 9500 28687 9503
rect 28902 9500 28908 9512
rect 28675 9472 28908 9500
rect 28675 9469 28687 9472
rect 28629 9463 28687 9469
rect 28902 9460 28908 9472
rect 28960 9460 28966 9512
rect 29086 9460 29092 9512
rect 29144 9500 29150 9512
rect 29273 9503 29331 9509
rect 29273 9500 29285 9503
rect 29144 9472 29285 9500
rect 29144 9460 29150 9472
rect 29273 9469 29285 9472
rect 29319 9469 29331 9503
rect 29273 9463 29331 9469
rect 4982 9392 4988 9444
rect 5040 9432 5046 9444
rect 25133 9435 25191 9441
rect 25133 9432 25145 9435
rect 5040 9404 25145 9432
rect 5040 9392 5046 9404
rect 25133 9401 25145 9404
rect 25179 9401 25191 9435
rect 25133 9395 25191 9401
rect 27430 9392 27436 9444
rect 27488 9432 27494 9444
rect 29380 9432 29408 9540
rect 30484 9540 32036 9568
rect 29914 9460 29920 9512
rect 29972 9509 29978 9512
rect 29972 9500 29983 9509
rect 30484 9500 30512 9540
rect 32030 9528 32036 9540
rect 32088 9528 32094 9580
rect 29972 9472 30512 9500
rect 30561 9503 30619 9509
rect 29972 9463 29983 9472
rect 30561 9469 30573 9503
rect 30607 9500 30619 9503
rect 31662 9500 31668 9512
rect 30607 9472 31668 9500
rect 30607 9469 30619 9472
rect 30561 9463 30619 9469
rect 29972 9460 29978 9463
rect 31662 9460 31668 9472
rect 31720 9460 31726 9512
rect 30466 9432 30472 9444
rect 27488 9404 29132 9432
rect 29380 9404 30472 9432
rect 27488 9392 27494 9404
rect 21266 9324 21272 9376
rect 21324 9364 21330 9376
rect 23845 9367 23903 9373
rect 23845 9364 23857 9367
rect 21324 9336 23857 9364
rect 21324 9324 21330 9336
rect 23845 9333 23857 9336
rect 23891 9333 23903 9367
rect 23845 9327 23903 9333
rect 25406 9324 25412 9376
rect 25464 9364 25470 9376
rect 26421 9367 26479 9373
rect 26421 9364 26433 9367
rect 25464 9336 26433 9364
rect 25464 9324 25470 9336
rect 26421 9333 26433 9336
rect 26467 9333 26479 9367
rect 26421 9327 26479 9333
rect 27246 9324 27252 9376
rect 27304 9364 27310 9376
rect 27801 9367 27859 9373
rect 27801 9364 27813 9367
rect 27304 9336 27813 9364
rect 27304 9324 27310 9336
rect 27801 9333 27813 9336
rect 27847 9333 27859 9367
rect 27801 9327 27859 9333
rect 28445 9367 28503 9373
rect 28445 9333 28457 9367
rect 28491 9364 28503 9367
rect 28534 9364 28540 9376
rect 28491 9336 28540 9364
rect 28491 9333 28503 9336
rect 28445 9327 28503 9333
rect 28534 9324 28540 9336
rect 28592 9324 28598 9376
rect 29104 9373 29132 9404
rect 30466 9392 30472 9404
rect 30524 9392 30530 9444
rect 29089 9367 29147 9373
rect 29089 9333 29101 9367
rect 29135 9333 29147 9367
rect 29089 9327 29147 9333
rect 29178 9324 29184 9376
rect 29236 9364 29242 9376
rect 29733 9367 29791 9373
rect 29733 9364 29745 9367
rect 29236 9336 29745 9364
rect 29236 9324 29242 9336
rect 29733 9333 29745 9336
rect 29779 9333 29791 9367
rect 29733 9327 29791 9333
rect 1104 9274 38824 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 38824 9274
rect 1104 9200 38824 9222
rect 22370 9120 22376 9172
rect 22428 9160 22434 9172
rect 22830 9160 22836 9172
rect 22428 9132 22836 9160
rect 22428 9120 22434 9132
rect 22830 9120 22836 9132
rect 22888 9120 22894 9172
rect 25424 9132 31340 9160
rect 25424 9104 25452 9132
rect 25406 9092 25412 9104
rect 23032 9064 25412 9092
rect 20714 8984 20720 9036
rect 20772 9024 20778 9036
rect 23032 9033 23060 9064
rect 25406 9052 25412 9064
rect 25464 9052 25470 9104
rect 26234 9052 26240 9104
rect 26292 9052 26298 9104
rect 26697 9095 26755 9101
rect 26697 9061 26709 9095
rect 26743 9092 26755 9095
rect 30282 9092 30288 9104
rect 26743 9064 30288 9092
rect 26743 9061 26755 9064
rect 26697 9055 26755 9061
rect 30282 9052 30288 9064
rect 30340 9052 30346 9104
rect 23017 9027 23075 9033
rect 23017 9024 23029 9027
rect 20772 8996 23029 9024
rect 20772 8984 20778 8996
rect 23017 8993 23029 8996
rect 23063 8993 23075 9027
rect 23658 9024 23664 9036
rect 23619 8996 23664 9024
rect 23017 8987 23075 8993
rect 23658 8984 23664 8996
rect 23716 8984 23722 9036
rect 24121 9027 24179 9033
rect 24121 8993 24133 9027
rect 24167 8993 24179 9027
rect 24121 8987 24179 8993
rect 27433 9027 27491 9033
rect 27433 8993 27445 9027
rect 27479 9024 27491 9027
rect 27614 9024 27620 9036
rect 27479 8996 27620 9024
rect 27479 8993 27491 8996
rect 27433 8987 27491 8993
rect 23842 8916 23848 8968
rect 23900 8956 23906 8968
rect 24136 8956 24164 8987
rect 27614 8984 27620 8996
rect 27672 8984 27678 9036
rect 28074 9024 28080 9036
rect 28035 8996 28080 9024
rect 28074 8984 28080 8996
rect 28132 8984 28138 9036
rect 28902 9024 28908 9036
rect 28863 8996 28908 9024
rect 28902 8984 28908 8996
rect 28960 8984 28966 9036
rect 29086 8984 29092 9036
rect 29144 9024 29150 9036
rect 29549 9027 29607 9033
rect 29549 9024 29561 9027
rect 29144 8996 29561 9024
rect 29144 8984 29150 8996
rect 29549 8993 29561 8996
rect 29595 9024 29607 9027
rect 30190 9024 30196 9036
rect 29595 8996 30196 9024
rect 29595 8993 29607 8996
rect 29549 8987 29607 8993
rect 30190 8984 30196 8996
rect 30248 8984 30254 9036
rect 30650 9024 30656 9036
rect 30611 8996 30656 9024
rect 30650 8984 30656 8996
rect 30708 8984 30714 9036
rect 31312 9033 31340 9132
rect 31297 9027 31355 9033
rect 31297 8993 31309 9027
rect 31343 9024 31355 9027
rect 37826 9024 37832 9036
rect 31343 8996 37832 9024
rect 31343 8993 31355 8996
rect 31297 8987 31355 8993
rect 37826 8984 37832 8996
rect 37884 8984 37890 9036
rect 26973 8959 27031 8965
rect 23900 8928 26924 8956
rect 23900 8916 23906 8928
rect 26896 8888 26924 8928
rect 26973 8925 26985 8959
rect 27019 8956 27031 8959
rect 27798 8956 27804 8968
rect 27019 8928 27804 8956
rect 27019 8925 27031 8928
rect 26973 8919 27031 8925
rect 27798 8916 27804 8928
rect 27856 8916 27862 8968
rect 27890 8916 27896 8968
rect 27948 8956 27954 8968
rect 30098 8956 30104 8968
rect 27948 8928 30104 8956
rect 27948 8916 27954 8928
rect 30098 8916 30104 8928
rect 30156 8956 30162 8968
rect 30668 8956 30696 8984
rect 31478 8956 31484 8968
rect 30156 8928 30604 8956
rect 30668 8928 31484 8956
rect 30156 8916 30162 8928
rect 27246 8888 27252 8900
rect 26896 8860 27252 8888
rect 27246 8848 27252 8860
rect 27304 8848 27310 8900
rect 28261 8891 28319 8897
rect 28261 8857 28273 8891
rect 28307 8888 28319 8891
rect 30466 8888 30472 8900
rect 28307 8860 30328 8888
rect 30427 8860 30472 8888
rect 28307 8857 28319 8860
rect 28261 8851 28319 8857
rect 23477 8823 23535 8829
rect 23477 8789 23489 8823
rect 23523 8820 23535 8823
rect 23658 8820 23664 8832
rect 23523 8792 23664 8820
rect 23523 8789 23535 8792
rect 23477 8783 23535 8789
rect 23658 8780 23664 8792
rect 23716 8780 23722 8832
rect 24305 8823 24363 8829
rect 24305 8789 24317 8823
rect 24351 8820 24363 8823
rect 24762 8820 24768 8832
rect 24351 8792 24768 8820
rect 24351 8789 24363 8792
rect 24305 8783 24363 8789
rect 24762 8780 24768 8792
rect 24820 8780 24826 8832
rect 25038 8780 25044 8832
rect 25096 8820 25102 8832
rect 25225 8823 25283 8829
rect 25225 8820 25237 8823
rect 25096 8792 25237 8820
rect 25096 8780 25102 8792
rect 25225 8789 25237 8792
rect 25271 8789 25283 8823
rect 25225 8783 25283 8789
rect 27617 8823 27675 8829
rect 27617 8789 27629 8823
rect 27663 8820 27675 8823
rect 28074 8820 28080 8832
rect 27663 8792 28080 8820
rect 27663 8789 27675 8792
rect 27617 8783 27675 8789
rect 28074 8780 28080 8792
rect 28132 8780 28138 8832
rect 28166 8780 28172 8832
rect 28224 8820 28230 8832
rect 28721 8823 28779 8829
rect 28721 8820 28733 8823
rect 28224 8792 28733 8820
rect 28224 8780 28230 8792
rect 28721 8789 28733 8792
rect 28767 8789 28779 8823
rect 28721 8783 28779 8789
rect 28902 8780 28908 8832
rect 28960 8820 28966 8832
rect 29365 8823 29423 8829
rect 29365 8820 29377 8823
rect 28960 8792 29377 8820
rect 28960 8780 28966 8792
rect 29365 8789 29377 8792
rect 29411 8789 29423 8823
rect 30300 8820 30328 8860
rect 30466 8848 30472 8860
rect 30524 8848 30530 8900
rect 30374 8820 30380 8832
rect 30300 8792 30380 8820
rect 29365 8783 29423 8789
rect 30374 8780 30380 8792
rect 30432 8780 30438 8832
rect 30576 8820 30604 8928
rect 31478 8916 31484 8928
rect 31536 8916 31542 8968
rect 30834 8848 30840 8900
rect 30892 8888 30898 8900
rect 31113 8891 31171 8897
rect 31113 8888 31125 8891
rect 30892 8860 31125 8888
rect 30892 8848 30898 8860
rect 31113 8857 31125 8860
rect 31159 8857 31171 8891
rect 31113 8851 31171 8857
rect 35434 8820 35440 8832
rect 30576 8792 35440 8820
rect 35434 8780 35440 8792
rect 35492 8780 35498 8832
rect 1104 8730 38824 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 38824 8730
rect 1104 8656 38824 8678
rect 27706 8576 27712 8628
rect 27764 8616 27770 8628
rect 27764 8588 29500 8616
rect 27764 8576 27770 8588
rect 20438 8508 20444 8560
rect 20496 8548 20502 8560
rect 24121 8551 24179 8557
rect 24121 8548 24133 8551
rect 20496 8520 24133 8548
rect 20496 8508 20502 8520
rect 24121 8517 24133 8520
rect 24167 8517 24179 8551
rect 24121 8511 24179 8517
rect 24302 8508 24308 8560
rect 24360 8548 24366 8560
rect 24360 8520 25176 8548
rect 24360 8508 24366 8520
rect 25148 8489 25176 8520
rect 25133 8483 25191 8489
rect 25133 8449 25145 8483
rect 25179 8449 25191 8483
rect 25133 8443 25191 8449
rect 26881 8483 26939 8489
rect 26881 8449 26893 8483
rect 26927 8480 26939 8483
rect 28810 8480 28816 8492
rect 26927 8452 28816 8480
rect 26927 8449 26939 8452
rect 26881 8443 26939 8449
rect 28810 8440 28816 8452
rect 28868 8440 28874 8492
rect 29178 8440 29184 8492
rect 29236 8480 29242 8492
rect 29273 8483 29331 8489
rect 29273 8480 29285 8483
rect 29236 8452 29285 8480
rect 29236 8440 29242 8452
rect 29273 8449 29285 8452
rect 29319 8449 29331 8483
rect 29472 8480 29500 8588
rect 30098 8576 30104 8628
rect 30156 8616 30162 8628
rect 30193 8619 30251 8625
rect 30193 8616 30205 8619
rect 30156 8588 30205 8616
rect 30156 8576 30162 8588
rect 30193 8585 30205 8588
rect 30239 8585 30251 8619
rect 30193 8579 30251 8585
rect 31202 8576 31208 8628
rect 31260 8616 31266 8628
rect 31297 8619 31355 8625
rect 31297 8616 31309 8619
rect 31260 8588 31309 8616
rect 31260 8576 31266 8588
rect 31297 8585 31309 8588
rect 31343 8585 31355 8619
rect 31849 8619 31907 8625
rect 31849 8616 31861 8619
rect 31297 8579 31355 8585
rect 31726 8588 31861 8616
rect 29546 8508 29552 8560
rect 29604 8548 29610 8560
rect 31726 8548 31754 8588
rect 31849 8585 31861 8588
rect 31895 8585 31907 8619
rect 31849 8579 31907 8585
rect 29604 8520 31754 8548
rect 29604 8508 29610 8520
rect 32674 8480 32680 8492
rect 29472 8452 32680 8480
rect 29273 8443 29331 8449
rect 22833 8415 22891 8421
rect 22833 8381 22845 8415
rect 22879 8412 22891 8415
rect 22922 8412 22928 8424
rect 22879 8384 22928 8412
rect 22879 8381 22891 8384
rect 22833 8375 22891 8381
rect 22922 8372 22928 8384
rect 22980 8372 22986 8424
rect 23661 8415 23719 8421
rect 23661 8381 23673 8415
rect 23707 8412 23719 8415
rect 23842 8412 23848 8424
rect 23707 8384 23848 8412
rect 23707 8381 23719 8384
rect 23661 8375 23719 8381
rect 22002 8304 22008 8356
rect 22060 8344 22066 8356
rect 23676 8344 23704 8375
rect 23842 8372 23848 8384
rect 23900 8372 23906 8424
rect 24305 8415 24363 8421
rect 24305 8381 24317 8415
rect 24351 8381 24363 8415
rect 24305 8375 24363 8381
rect 22060 8316 23704 8344
rect 22060 8304 22066 8316
rect 23014 8276 23020 8288
rect 22975 8248 23020 8276
rect 23014 8236 23020 8248
rect 23072 8236 23078 8288
rect 23474 8276 23480 8288
rect 23435 8248 23480 8276
rect 23474 8236 23480 8248
rect 23532 8236 23538 8288
rect 24320 8276 24348 8375
rect 29546 8372 29552 8424
rect 29604 8412 29610 8424
rect 30024 8421 30052 8452
rect 32674 8440 32680 8452
rect 32732 8440 32738 8492
rect 30009 8415 30067 8421
rect 29604 8384 29649 8412
rect 29604 8372 29610 8384
rect 30009 8381 30021 8415
rect 30055 8381 30067 8415
rect 31386 8412 31392 8424
rect 31347 8384 31392 8412
rect 30009 8375 30067 8381
rect 31386 8372 31392 8384
rect 31444 8372 31450 8424
rect 31662 8372 31668 8424
rect 31720 8412 31726 8424
rect 32033 8415 32091 8421
rect 32033 8412 32045 8415
rect 31720 8384 32045 8412
rect 31720 8372 31726 8384
rect 32033 8381 32045 8384
rect 32079 8381 32091 8415
rect 32033 8375 32091 8381
rect 24394 8304 24400 8356
rect 24452 8344 24458 8356
rect 25409 8347 25467 8353
rect 25409 8344 25421 8347
rect 24452 8316 25421 8344
rect 24452 8304 24458 8316
rect 25409 8313 25421 8316
rect 25455 8313 25467 8347
rect 27890 8344 27896 8356
rect 26634 8316 27896 8344
rect 25409 8307 25467 8313
rect 27890 8304 27896 8316
rect 27948 8304 27954 8356
rect 35710 8344 35716 8356
rect 28842 8316 29224 8344
rect 24670 8276 24676 8288
rect 24320 8248 24676 8276
rect 24670 8236 24676 8248
rect 24728 8276 24734 8288
rect 25222 8276 25228 8288
rect 24728 8248 25228 8276
rect 24728 8236 24734 8248
rect 25222 8236 25228 8248
rect 25280 8236 25286 8288
rect 27798 8276 27804 8288
rect 27759 8248 27804 8276
rect 27798 8236 27804 8248
rect 27856 8236 27862 8288
rect 29196 8276 29224 8316
rect 29380 8316 35716 8344
rect 29380 8276 29408 8316
rect 35710 8304 35716 8316
rect 35768 8304 35774 8356
rect 29196 8248 29408 8276
rect 31478 8236 31484 8288
rect 31536 8276 31542 8288
rect 33134 8276 33140 8288
rect 31536 8248 33140 8276
rect 31536 8236 31542 8248
rect 33134 8236 33140 8248
rect 33192 8236 33198 8288
rect 1104 8186 38824 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 38824 8186
rect 1104 8112 38824 8134
rect 18966 8032 18972 8084
rect 19024 8072 19030 8084
rect 22557 8075 22615 8081
rect 22557 8072 22569 8075
rect 19024 8044 22569 8072
rect 19024 8032 19030 8044
rect 22557 8041 22569 8044
rect 22603 8041 22615 8075
rect 36538 8072 36544 8084
rect 22557 8035 22615 8041
rect 26712 8044 36544 8072
rect 19426 7964 19432 8016
rect 19484 8004 19490 8016
rect 19484 7976 22784 8004
rect 19484 7964 19490 7976
rect 21277 7939 21335 7945
rect 21277 7905 21289 7939
rect 21323 7936 21335 7939
rect 21323 7908 21496 7936
rect 21323 7905 21335 7908
rect 21277 7899 21335 7905
rect 21468 7868 21496 7908
rect 21542 7896 21548 7948
rect 21600 7936 21606 7948
rect 22097 7939 22155 7945
rect 22097 7936 22109 7939
rect 21600 7908 22109 7936
rect 21600 7896 21606 7908
rect 22097 7905 22109 7908
rect 22143 7936 22155 7939
rect 22143 7908 22600 7936
rect 22143 7905 22155 7908
rect 22097 7899 22155 7905
rect 22370 7868 22376 7880
rect 21468 7840 22376 7868
rect 22370 7828 22376 7840
rect 22428 7828 22434 7880
rect 21453 7803 21511 7809
rect 21453 7769 21465 7803
rect 21499 7800 21511 7803
rect 22462 7800 22468 7812
rect 21499 7772 22468 7800
rect 21499 7769 21511 7772
rect 21453 7763 21511 7769
rect 22462 7760 22468 7772
rect 22520 7760 22526 7812
rect 18230 7692 18236 7744
rect 18288 7732 18294 7744
rect 21542 7732 21548 7744
rect 18288 7704 21548 7732
rect 18288 7692 18294 7704
rect 21542 7692 21548 7704
rect 21600 7692 21606 7744
rect 21910 7732 21916 7744
rect 21871 7704 21916 7732
rect 21910 7692 21916 7704
rect 21968 7692 21974 7744
rect 22572 7732 22600 7908
rect 22756 7868 22784 7976
rect 23014 7964 23020 8016
rect 23072 7964 23078 8016
rect 26712 7990 26740 8044
rect 36538 8032 36544 8044
rect 36596 8032 36602 8084
rect 27798 7964 27804 8016
rect 27856 8004 27862 8016
rect 28077 8007 28135 8013
rect 28077 8004 28089 8007
rect 27856 7976 28089 8004
rect 27856 7964 27862 7976
rect 28077 7973 28089 7976
rect 28123 7973 28135 8007
rect 28077 7967 28135 7973
rect 28626 7964 28632 8016
rect 28684 7964 28690 8016
rect 32490 8004 32496 8016
rect 29564 7976 32496 8004
rect 24302 7896 24308 7948
rect 24360 7936 24366 7948
rect 24360 7908 24405 7936
rect 24360 7896 24366 7908
rect 24029 7871 24087 7877
rect 24029 7868 24041 7871
rect 22756 7840 24041 7868
rect 24029 7837 24041 7840
rect 24075 7837 24087 7871
rect 24029 7831 24087 7837
rect 25225 7871 25283 7877
rect 25225 7837 25237 7871
rect 25271 7837 25283 7871
rect 25498 7868 25504 7880
rect 25459 7840 25504 7868
rect 25225 7831 25283 7837
rect 23566 7732 23572 7744
rect 22572 7704 23572 7732
rect 23566 7692 23572 7704
rect 23624 7692 23630 7744
rect 25240 7732 25268 7831
rect 25498 7828 25504 7840
rect 25556 7828 25562 7880
rect 27706 7828 27712 7880
rect 27764 7868 27770 7880
rect 27801 7871 27859 7877
rect 27801 7868 27813 7871
rect 27764 7840 27813 7868
rect 27764 7828 27770 7840
rect 27801 7837 27813 7840
rect 27847 7837 27859 7871
rect 27801 7831 27859 7837
rect 28074 7828 28080 7880
rect 28132 7868 28138 7880
rect 29564 7877 29592 7976
rect 32490 7964 32496 7976
rect 32548 7964 32554 8016
rect 30650 7936 30656 7948
rect 30611 7908 30656 7936
rect 30650 7896 30656 7908
rect 30708 7896 30714 7948
rect 31289 7939 31347 7945
rect 31289 7905 31301 7939
rect 31335 7905 31347 7939
rect 31289 7899 31347 7905
rect 31941 7939 31999 7945
rect 31941 7905 31953 7939
rect 31987 7936 31999 7939
rect 32030 7936 32036 7948
rect 31987 7908 32036 7936
rect 31987 7905 31999 7908
rect 31941 7899 31999 7905
rect 29549 7871 29607 7877
rect 28132 7840 29132 7868
rect 28132 7828 28138 7840
rect 27724 7800 27752 7828
rect 26528 7772 27752 7800
rect 29104 7800 29132 7840
rect 29549 7837 29561 7871
rect 29595 7837 29607 7871
rect 29549 7831 29607 7837
rect 30190 7828 30196 7880
rect 30248 7868 30254 7880
rect 31312 7868 31340 7899
rect 32030 7896 32036 7908
rect 32088 7896 32094 7948
rect 32585 7939 32643 7945
rect 32585 7905 32597 7939
rect 32631 7936 32643 7939
rect 33134 7936 33140 7948
rect 32631 7908 33140 7936
rect 32631 7905 32643 7908
rect 32585 7899 32643 7905
rect 33134 7896 33140 7908
rect 33192 7896 33198 7948
rect 33229 7939 33287 7945
rect 33229 7905 33241 7939
rect 33275 7936 33287 7939
rect 34606 7936 34612 7948
rect 33275 7908 34612 7936
rect 33275 7905 33287 7908
rect 33229 7899 33287 7905
rect 34606 7896 34612 7908
rect 34664 7896 34670 7948
rect 30248 7840 31340 7868
rect 30248 7828 30254 7840
rect 31570 7828 31576 7880
rect 31628 7868 31634 7880
rect 31628 7840 33088 7868
rect 31628 7828 31634 7840
rect 30834 7800 30840 7812
rect 29104 7772 30840 7800
rect 26528 7732 26556 7772
rect 30834 7760 30840 7772
rect 30892 7760 30898 7812
rect 30926 7760 30932 7812
rect 30984 7800 30990 7812
rect 33060 7809 33088 7840
rect 31757 7803 31815 7809
rect 31757 7800 31769 7803
rect 30984 7772 31769 7800
rect 30984 7760 30990 7772
rect 31757 7769 31769 7772
rect 31803 7769 31815 7803
rect 31757 7763 31815 7769
rect 33045 7803 33103 7809
rect 33045 7769 33057 7803
rect 33091 7769 33103 7803
rect 33045 7763 33103 7769
rect 26970 7732 26976 7744
rect 25240 7704 26556 7732
rect 26931 7704 26976 7732
rect 26970 7692 26976 7704
rect 27028 7692 27034 7744
rect 27890 7692 27896 7744
rect 27948 7732 27954 7744
rect 30469 7735 30527 7741
rect 30469 7732 30481 7735
rect 27948 7704 30481 7732
rect 27948 7692 27954 7704
rect 30469 7701 30481 7704
rect 30515 7701 30527 7735
rect 31110 7732 31116 7744
rect 31071 7704 31116 7732
rect 30469 7695 30527 7701
rect 31110 7692 31116 7704
rect 31168 7692 31174 7744
rect 31846 7692 31852 7744
rect 31904 7732 31910 7744
rect 32401 7735 32459 7741
rect 32401 7732 32413 7735
rect 31904 7704 32413 7732
rect 31904 7692 31910 7704
rect 32401 7701 32413 7704
rect 32447 7701 32459 7735
rect 32401 7695 32459 7701
rect 1104 7642 38824 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 38824 7642
rect 1104 7568 38824 7590
rect 20901 7531 20959 7537
rect 20901 7497 20913 7531
rect 20947 7528 20959 7531
rect 25406 7528 25412 7540
rect 20947 7500 25412 7528
rect 20947 7497 20959 7500
rect 20901 7491 20959 7497
rect 21450 7420 21456 7472
rect 21508 7460 21514 7472
rect 23569 7463 23627 7469
rect 23569 7460 23581 7463
rect 21508 7432 23581 7460
rect 21508 7420 21514 7432
rect 23569 7429 23581 7432
rect 23615 7429 23627 7463
rect 23569 7423 23627 7429
rect 17862 7352 17868 7404
rect 17920 7392 17926 7404
rect 23109 7395 23167 7401
rect 23109 7392 23121 7395
rect 17920 7364 23121 7392
rect 17920 7352 17926 7364
rect 23109 7361 23121 7364
rect 23155 7361 23167 7395
rect 23676 7392 23704 7500
rect 25406 7488 25412 7500
rect 25464 7488 25470 7540
rect 26234 7488 26240 7540
rect 26292 7528 26298 7540
rect 30653 7531 30711 7537
rect 30653 7528 30665 7531
rect 26292 7500 30665 7528
rect 26292 7488 26298 7500
rect 30653 7497 30665 7500
rect 30699 7497 30711 7531
rect 30653 7491 30711 7497
rect 30742 7488 30748 7540
rect 30800 7528 30806 7540
rect 31941 7531 31999 7537
rect 31941 7528 31953 7531
rect 30800 7500 31953 7528
rect 30800 7488 30806 7500
rect 31941 7497 31953 7500
rect 31987 7497 31999 7531
rect 31941 7491 31999 7497
rect 29914 7420 29920 7472
rect 29972 7460 29978 7472
rect 30926 7460 30932 7472
rect 29972 7432 30932 7460
rect 29972 7420 29978 7432
rect 30926 7420 30932 7432
rect 30984 7420 30990 7472
rect 23109 7355 23167 7361
rect 23400 7364 23704 7392
rect 20257 7327 20315 7333
rect 20257 7293 20269 7327
rect 20303 7324 20315 7327
rect 20622 7324 20628 7336
rect 20303 7296 20628 7324
rect 20303 7293 20315 7296
rect 20257 7287 20315 7293
rect 20622 7284 20628 7296
rect 20680 7284 20686 7336
rect 20833 7327 20891 7333
rect 20833 7293 20845 7327
rect 20879 7324 20891 7327
rect 21358 7324 21364 7336
rect 20879 7296 21364 7324
rect 20879 7293 20891 7296
rect 20833 7287 20891 7293
rect 21358 7284 21364 7296
rect 21416 7284 21422 7336
rect 21453 7327 21511 7333
rect 21453 7293 21465 7327
rect 21499 7324 21511 7327
rect 22094 7324 22100 7336
rect 21499 7296 22100 7324
rect 21499 7293 21511 7296
rect 21453 7287 21511 7293
rect 22094 7284 22100 7296
rect 22152 7324 22158 7336
rect 22922 7324 22928 7336
rect 22152 7296 22928 7324
rect 22152 7284 22158 7296
rect 22922 7284 22928 7296
rect 22980 7284 22986 7336
rect 23014 7284 23020 7336
rect 23072 7324 23078 7336
rect 23400 7333 23428 7364
rect 24302 7352 24308 7404
rect 24360 7392 24366 7404
rect 24578 7392 24584 7404
rect 24360 7364 24584 7392
rect 24360 7352 24366 7364
rect 24578 7352 24584 7364
rect 24636 7352 24642 7404
rect 28626 7352 28632 7404
rect 28684 7392 28690 7404
rect 28684 7364 30052 7392
rect 28684 7352 28690 7364
rect 23293 7327 23351 7333
rect 23293 7324 23305 7327
rect 23072 7296 23305 7324
rect 23072 7284 23078 7296
rect 23293 7293 23305 7296
rect 23339 7293 23351 7327
rect 23293 7287 23351 7293
rect 23385 7327 23443 7333
rect 23385 7293 23397 7327
rect 23431 7293 23443 7327
rect 23385 7287 23443 7293
rect 23661 7327 23719 7333
rect 23661 7293 23673 7327
rect 23707 7324 23719 7327
rect 23934 7324 23940 7336
rect 23707 7296 23940 7324
rect 23707 7293 23719 7296
rect 23661 7287 23719 7293
rect 23934 7284 23940 7296
rect 23992 7284 23998 7336
rect 29546 7284 29552 7336
rect 29604 7324 29610 7336
rect 30024 7333 30052 7364
rect 30190 7352 30196 7404
rect 30248 7392 30254 7404
rect 36906 7392 36912 7404
rect 30248 7364 36912 7392
rect 30248 7352 30254 7364
rect 30009 7327 30067 7333
rect 29604 7296 29649 7324
rect 29604 7284 29610 7296
rect 30009 7293 30021 7327
rect 30055 7293 30067 7327
rect 30834 7324 30840 7336
rect 30747 7296 30840 7324
rect 30009 7287 30067 7293
rect 30834 7284 30840 7296
rect 30892 7284 30898 7336
rect 30926 7284 30932 7336
rect 30984 7324 30990 7336
rect 31386 7324 31392 7336
rect 30984 7296 31392 7324
rect 30984 7284 30990 7296
rect 31386 7284 31392 7296
rect 31444 7324 31450 7336
rect 32140 7333 32168 7364
rect 36906 7352 36912 7364
rect 36964 7352 36970 7404
rect 31481 7327 31539 7333
rect 31481 7324 31493 7327
rect 31444 7296 31493 7324
rect 31444 7284 31450 7296
rect 31481 7293 31493 7296
rect 31527 7293 31539 7327
rect 31481 7287 31539 7293
rect 32125 7327 32183 7333
rect 32125 7293 32137 7327
rect 32171 7293 32183 7327
rect 32125 7287 32183 7293
rect 33134 7284 33140 7336
rect 33192 7324 33198 7336
rect 33229 7327 33287 7333
rect 33229 7324 33241 7327
rect 33192 7296 33241 7324
rect 33192 7284 33198 7296
rect 33229 7293 33241 7296
rect 33275 7293 33287 7327
rect 33229 7287 33287 7293
rect 16022 7216 16028 7268
rect 16080 7256 16086 7268
rect 24854 7256 24860 7268
rect 16080 7228 23704 7256
rect 24815 7228 24860 7256
rect 16080 7216 16086 7228
rect 20070 7188 20076 7200
rect 20031 7160 20076 7188
rect 20070 7148 20076 7160
rect 20128 7148 20134 7200
rect 21637 7191 21695 7197
rect 21637 7157 21649 7191
rect 21683 7188 21695 7191
rect 21818 7188 21824 7200
rect 21683 7160 21824 7188
rect 21683 7157 21695 7160
rect 21637 7151 21695 7157
rect 21818 7148 21824 7160
rect 21876 7148 21882 7200
rect 23676 7188 23704 7228
rect 24854 7216 24860 7228
rect 24912 7216 24918 7268
rect 25332 7188 25360 7242
rect 28534 7216 28540 7268
rect 28592 7216 28598 7268
rect 29273 7259 29331 7265
rect 29273 7225 29285 7259
rect 29319 7225 29331 7259
rect 30852 7256 30880 7284
rect 32950 7256 32956 7268
rect 30852 7228 32956 7256
rect 29273 7219 29331 7225
rect 23676 7160 25360 7188
rect 25774 7148 25780 7200
rect 25832 7188 25838 7200
rect 26329 7191 26387 7197
rect 26329 7188 26341 7191
rect 25832 7160 26341 7188
rect 25832 7148 25838 7160
rect 26329 7157 26341 7160
rect 26375 7157 26387 7191
rect 26329 7151 26387 7157
rect 26418 7148 26424 7200
rect 26476 7188 26482 7200
rect 27801 7191 27859 7197
rect 27801 7188 27813 7191
rect 26476 7160 27813 7188
rect 26476 7148 26482 7160
rect 27801 7157 27813 7160
rect 27847 7157 27859 7191
rect 27801 7151 27859 7157
rect 27890 7148 27896 7200
rect 27948 7188 27954 7200
rect 29288 7188 29316 7219
rect 32950 7216 32956 7228
rect 33008 7216 33014 7268
rect 33244 7256 33272 7287
rect 33686 7284 33692 7336
rect 33744 7324 33750 7336
rect 33873 7327 33931 7333
rect 33873 7324 33885 7327
rect 33744 7296 33885 7324
rect 33744 7284 33750 7296
rect 33873 7293 33885 7296
rect 33919 7293 33931 7327
rect 33873 7287 33931 7293
rect 34146 7256 34152 7268
rect 33244 7228 34152 7256
rect 34146 7216 34152 7228
rect 34204 7216 34210 7268
rect 30190 7188 30196 7200
rect 27948 7160 29316 7188
rect 30151 7160 30196 7188
rect 27948 7148 27954 7160
rect 30190 7148 30196 7160
rect 30248 7148 30254 7200
rect 30650 7148 30656 7200
rect 30708 7188 30714 7200
rect 30926 7188 30932 7200
rect 30708 7160 30932 7188
rect 30708 7148 30714 7160
rect 30926 7148 30932 7160
rect 30984 7148 30990 7200
rect 31294 7188 31300 7200
rect 31255 7160 31300 7188
rect 31294 7148 31300 7160
rect 31352 7148 31358 7200
rect 31938 7148 31944 7200
rect 31996 7188 32002 7200
rect 33045 7191 33103 7197
rect 33045 7188 33057 7191
rect 31996 7160 33057 7188
rect 31996 7148 32002 7160
rect 33045 7157 33057 7160
rect 33091 7157 33103 7191
rect 33045 7151 33103 7157
rect 33781 7191 33839 7197
rect 33781 7157 33793 7191
rect 33827 7188 33839 7191
rect 34054 7188 34060 7200
rect 33827 7160 34060 7188
rect 33827 7157 33839 7160
rect 33781 7151 33839 7157
rect 34054 7148 34060 7160
rect 34112 7148 34118 7200
rect 1104 7098 38824 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 38824 7098
rect 1104 7024 38824 7046
rect 28166 6984 28172 6996
rect 24044 6956 28172 6984
rect 23106 6916 23112 6928
rect 21850 6888 23112 6916
rect 23106 6876 23112 6888
rect 23164 6876 23170 6928
rect 24044 6902 24072 6956
rect 28166 6944 28172 6956
rect 28224 6944 28230 6996
rect 30006 6944 30012 6996
rect 30064 6984 30070 6996
rect 31570 6984 31576 6996
rect 30064 6956 31576 6984
rect 30064 6944 30070 6956
rect 31570 6944 31576 6956
rect 31628 6944 31634 6996
rect 32030 6944 32036 6996
rect 32088 6984 32094 6996
rect 33505 6987 33563 6993
rect 33505 6984 33517 6987
rect 32088 6956 33517 6984
rect 32088 6944 32094 6956
rect 33505 6953 33517 6956
rect 33551 6984 33563 6987
rect 34698 6984 34704 6996
rect 33551 6956 34704 6984
rect 33551 6953 33563 6956
rect 33505 6947 33563 6953
rect 34698 6944 34704 6956
rect 34756 6944 34762 6996
rect 26418 6916 26424 6928
rect 24136 6888 26424 6916
rect 19886 6740 19892 6792
rect 19944 6780 19950 6792
rect 20349 6783 20407 6789
rect 20349 6780 20361 6783
rect 19944 6752 20361 6780
rect 19944 6740 19950 6752
rect 20349 6749 20361 6752
rect 20395 6749 20407 6783
rect 20625 6783 20683 6789
rect 20625 6780 20637 6783
rect 20349 6743 20407 6749
rect 20456 6752 20637 6780
rect 16482 6672 16488 6724
rect 16540 6712 16546 6724
rect 20456 6712 20484 6752
rect 20625 6749 20637 6752
rect 20671 6749 20683 6783
rect 22554 6780 22560 6792
rect 22515 6752 22560 6780
rect 20625 6743 20683 6749
rect 22554 6740 22560 6752
rect 22612 6740 22618 6792
rect 22833 6783 22891 6789
rect 22833 6749 22845 6783
rect 22879 6780 22891 6783
rect 24136 6780 24164 6888
rect 26418 6876 26424 6888
rect 26476 6876 26482 6928
rect 28902 6916 28908 6928
rect 27370 6888 28908 6916
rect 28902 6876 28908 6888
rect 28960 6876 28966 6928
rect 30190 6876 30196 6928
rect 30248 6916 30254 6928
rect 30248 6888 30774 6916
rect 30248 6876 30254 6888
rect 31662 6876 31668 6928
rect 31720 6916 31726 6928
rect 31720 6888 33456 6916
rect 31720 6876 31726 6888
rect 33428 6860 33456 6888
rect 24210 6808 24216 6860
rect 24268 6848 24274 6860
rect 25685 6851 25743 6857
rect 25685 6848 25697 6851
rect 24268 6820 25697 6848
rect 24268 6808 24274 6820
rect 25685 6817 25697 6820
rect 25731 6848 25743 6851
rect 25731 6820 26648 6848
rect 25731 6817 25743 6820
rect 25685 6811 25743 6817
rect 22879 6752 24164 6780
rect 24305 6783 24363 6789
rect 22879 6749 22891 6752
rect 22833 6743 22891 6749
rect 24305 6749 24317 6783
rect 24351 6780 24363 6783
rect 24394 6780 24400 6792
rect 24351 6752 24400 6780
rect 24351 6749 24363 6752
rect 24305 6743 24363 6749
rect 24394 6740 24400 6752
rect 24452 6740 24458 6792
rect 25593 6783 25651 6789
rect 25593 6749 25605 6783
rect 25639 6780 25651 6783
rect 26329 6783 26387 6789
rect 26329 6780 26341 6783
rect 25639 6752 26341 6780
rect 25639 6749 25651 6752
rect 25593 6743 25651 6749
rect 26329 6749 26341 6752
rect 26375 6749 26387 6783
rect 26620 6780 26648 6820
rect 28534 6808 28540 6860
rect 28592 6848 28598 6860
rect 28629 6851 28687 6857
rect 28629 6848 28641 6851
rect 28592 6820 28641 6848
rect 28592 6808 28598 6820
rect 28629 6817 28641 6820
rect 28675 6848 28687 6851
rect 29273 6851 29331 6857
rect 29273 6848 29285 6851
rect 28675 6820 29285 6848
rect 28675 6817 28687 6820
rect 28629 6811 28687 6817
rect 29273 6817 29285 6820
rect 29319 6817 29331 6851
rect 29546 6848 29552 6860
rect 29273 6811 29331 6817
rect 29380 6820 29552 6848
rect 27338 6780 27344 6792
rect 26620 6752 27344 6780
rect 26329 6743 26387 6749
rect 27338 6740 27344 6752
rect 27396 6740 27402 6792
rect 27798 6780 27804 6792
rect 27759 6752 27804 6780
rect 27798 6740 27804 6752
rect 27856 6740 27862 6792
rect 28077 6783 28135 6789
rect 28077 6780 28089 6783
rect 28000 6752 28089 6780
rect 16540 6684 20484 6712
rect 16540 6672 16546 6684
rect 25222 6672 25228 6724
rect 25280 6712 25286 6724
rect 25869 6715 25927 6721
rect 25869 6712 25881 6715
rect 25280 6684 25881 6712
rect 25280 6672 25286 6684
rect 25869 6681 25881 6684
rect 25915 6681 25927 6715
rect 25869 6675 25927 6681
rect 22097 6647 22155 6653
rect 22097 6613 22109 6647
rect 22143 6644 22155 6647
rect 22186 6644 22192 6656
rect 22143 6616 22192 6644
rect 22143 6613 22155 6616
rect 22097 6607 22155 6613
rect 22186 6604 22192 6616
rect 22244 6604 22250 6656
rect 22922 6604 22928 6656
rect 22980 6644 22986 6656
rect 25593 6647 25651 6653
rect 25593 6644 25605 6647
rect 22980 6616 25605 6644
rect 22980 6604 22986 6616
rect 25593 6613 25605 6616
rect 25639 6613 25651 6647
rect 25593 6607 25651 6613
rect 27338 6604 27344 6656
rect 27396 6644 27402 6656
rect 27614 6644 27620 6656
rect 27396 6616 27620 6644
rect 27396 6604 27402 6616
rect 27614 6604 27620 6616
rect 27672 6604 27678 6656
rect 27706 6604 27712 6656
rect 27764 6644 27770 6656
rect 28000 6644 28028 6752
rect 28077 6749 28089 6752
rect 28123 6780 28135 6783
rect 29380 6780 29408 6820
rect 29546 6808 29552 6820
rect 29604 6808 29610 6860
rect 32306 6808 32312 6860
rect 32364 6848 32370 6860
rect 32674 6848 32680 6860
rect 32364 6820 32536 6848
rect 32635 6820 32680 6848
rect 32364 6808 32370 6820
rect 31478 6780 31484 6792
rect 28123 6752 29408 6780
rect 29472 6752 31484 6780
rect 28123 6749 28135 6752
rect 28077 6743 28135 6749
rect 29472 6721 29500 6752
rect 31478 6740 31484 6752
rect 31536 6740 31542 6792
rect 31570 6740 31576 6792
rect 31628 6780 31634 6792
rect 31846 6780 31852 6792
rect 31628 6752 31852 6780
rect 31628 6740 31634 6752
rect 31846 6740 31852 6752
rect 31904 6740 31910 6792
rect 32217 6783 32275 6789
rect 32217 6749 32229 6783
rect 32263 6780 32275 6783
rect 32398 6780 32404 6792
rect 32263 6752 32404 6780
rect 32263 6749 32275 6752
rect 32217 6743 32275 6749
rect 32398 6740 32404 6752
rect 32456 6740 32462 6792
rect 32508 6780 32536 6820
rect 32674 6808 32680 6820
rect 32732 6848 32738 6860
rect 33042 6848 33048 6860
rect 32732 6820 33048 6848
rect 32732 6808 32738 6820
rect 33042 6808 33048 6820
rect 33100 6848 33106 6860
rect 33321 6851 33379 6857
rect 33321 6848 33333 6851
rect 33100 6820 33333 6848
rect 33100 6808 33106 6820
rect 33321 6817 33333 6820
rect 33367 6817 33379 6851
rect 33321 6811 33379 6817
rect 33410 6808 33416 6860
rect 33468 6808 33474 6860
rect 34146 6848 34152 6860
rect 34107 6820 34152 6848
rect 34146 6808 34152 6820
rect 34204 6808 34210 6860
rect 34606 6848 34612 6860
rect 34519 6820 34612 6848
rect 34606 6808 34612 6820
rect 34664 6848 34670 6860
rect 35802 6848 35808 6860
rect 34664 6820 35808 6848
rect 34664 6808 34670 6820
rect 35802 6808 35808 6820
rect 35860 6808 35866 6860
rect 35894 6780 35900 6792
rect 32508 6752 35900 6780
rect 35894 6740 35900 6752
rect 35952 6740 35958 6792
rect 29457 6715 29515 6721
rect 29457 6681 29469 6715
rect 29503 6681 29515 6715
rect 29457 6675 29515 6681
rect 33134 6672 33140 6724
rect 33192 6712 33198 6724
rect 33965 6715 34023 6721
rect 33965 6712 33977 6715
rect 33192 6684 33977 6712
rect 33192 6672 33198 6684
rect 33965 6681 33977 6684
rect 34011 6681 34023 6715
rect 33965 6675 34023 6681
rect 27764 6616 28028 6644
rect 28813 6647 28871 6653
rect 27764 6604 27770 6616
rect 28813 6613 28825 6647
rect 28859 6644 28871 6647
rect 29270 6644 29276 6656
rect 28859 6616 29276 6644
rect 28859 6613 28871 6616
rect 28813 6607 28871 6613
rect 29270 6604 29276 6616
rect 29328 6604 29334 6656
rect 30469 6647 30527 6653
rect 30469 6613 30481 6647
rect 30515 6644 30527 6647
rect 30650 6644 30656 6656
rect 30515 6616 30656 6644
rect 30515 6613 30527 6616
rect 30469 6607 30527 6613
rect 30650 6604 30656 6616
rect 30708 6604 30714 6656
rect 31754 6604 31760 6656
rect 31812 6644 31818 6656
rect 31953 6647 32011 6653
rect 31953 6644 31965 6647
rect 31812 6616 31965 6644
rect 31812 6604 31818 6616
rect 31953 6613 31965 6616
rect 31999 6613 32011 6647
rect 31953 6607 32011 6613
rect 32766 6604 32772 6656
rect 32824 6644 32830 6656
rect 32861 6647 32919 6653
rect 32861 6644 32873 6647
rect 32824 6616 32873 6644
rect 32824 6604 32830 6616
rect 32861 6613 32873 6616
rect 32907 6613 32919 6647
rect 32861 6607 32919 6613
rect 34606 6604 34612 6656
rect 34664 6644 34670 6656
rect 34793 6647 34851 6653
rect 34793 6644 34805 6647
rect 34664 6616 34805 6644
rect 34664 6604 34670 6616
rect 34793 6613 34805 6616
rect 34839 6613 34851 6647
rect 34793 6607 34851 6613
rect 1104 6554 38824 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 38824 6554
rect 1104 6480 38824 6502
rect 20254 6400 20260 6452
rect 20312 6440 20318 6452
rect 22370 6440 22376 6452
rect 20312 6412 22376 6440
rect 20312 6400 20318 6412
rect 22370 6400 22376 6412
rect 22428 6400 22434 6452
rect 24673 6443 24731 6449
rect 22480 6412 24624 6440
rect 22094 6304 22100 6316
rect 19444 6276 22100 6304
rect 18874 6196 18880 6248
rect 18932 6236 18938 6248
rect 19444 6245 19472 6276
rect 22094 6264 22100 6276
rect 22152 6264 22158 6316
rect 19429 6239 19487 6245
rect 19429 6236 19441 6239
rect 18932 6208 19441 6236
rect 18932 6196 18938 6208
rect 19429 6205 19441 6208
rect 19475 6205 19487 6239
rect 19886 6236 19892 6248
rect 19847 6208 19892 6236
rect 19429 6199 19487 6205
rect 19886 6196 19892 6208
rect 19944 6196 19950 6248
rect 22480 6236 22508 6412
rect 24486 6372 24492 6384
rect 24228 6344 24492 6372
rect 22554 6264 22560 6316
rect 22612 6304 22618 6316
rect 22925 6307 22983 6313
rect 22925 6304 22937 6307
rect 22612 6276 22937 6304
rect 22612 6264 22618 6276
rect 22925 6273 22937 6276
rect 22971 6304 22983 6307
rect 24228 6304 24256 6344
rect 24486 6332 24492 6344
rect 24544 6332 24550 6384
rect 24596 6372 24624 6412
rect 24673 6409 24685 6443
rect 24719 6440 24731 6443
rect 25498 6440 25504 6452
rect 24719 6412 25504 6440
rect 24719 6409 24731 6412
rect 24673 6403 24731 6409
rect 25498 6400 25504 6412
rect 25556 6400 25562 6452
rect 27816 6412 31754 6440
rect 24946 6372 24952 6384
rect 24596 6344 24952 6372
rect 24946 6332 24952 6344
rect 25004 6332 25010 6384
rect 26881 6375 26939 6381
rect 26881 6341 26893 6375
rect 26927 6372 26939 6375
rect 27614 6372 27620 6384
rect 26927 6344 27620 6372
rect 26927 6341 26939 6344
rect 26881 6335 26939 6341
rect 27614 6332 27620 6344
rect 27672 6332 27678 6384
rect 27816 6304 27844 6412
rect 30009 6375 30067 6381
rect 30009 6341 30021 6375
rect 30055 6372 30067 6375
rect 30466 6372 30472 6384
rect 30055 6344 30472 6372
rect 30055 6341 30067 6344
rect 30009 6335 30067 6341
rect 30466 6332 30472 6344
rect 30524 6332 30530 6384
rect 31726 6372 31754 6412
rect 31846 6400 31852 6452
rect 31904 6440 31910 6452
rect 32214 6440 32220 6452
rect 31904 6412 32220 6440
rect 31904 6400 31910 6412
rect 32214 6400 32220 6412
rect 32272 6400 32278 6452
rect 32306 6400 32312 6452
rect 32364 6440 32370 6452
rect 34333 6443 34391 6449
rect 34333 6440 34345 6443
rect 32364 6412 34345 6440
rect 32364 6400 32370 6412
rect 34333 6409 34345 6412
rect 34379 6409 34391 6443
rect 34333 6403 34391 6409
rect 31726 6344 31984 6372
rect 22971 6276 24256 6304
rect 24320 6276 27844 6304
rect 22971 6273 22983 6276
rect 22925 6267 22983 6273
rect 21298 6208 22508 6236
rect 24320 6222 24348 6276
rect 28074 6264 28080 6316
rect 28132 6304 28138 6316
rect 29454 6304 29460 6316
rect 28132 6276 29460 6304
rect 28132 6264 28138 6276
rect 29454 6264 29460 6276
rect 29512 6264 29518 6316
rect 29549 6307 29607 6313
rect 29549 6273 29561 6307
rect 29595 6304 29607 6307
rect 30742 6304 30748 6316
rect 29595 6276 30748 6304
rect 29595 6273 29607 6276
rect 29549 6267 29607 6273
rect 30742 6264 30748 6276
rect 30800 6264 30806 6316
rect 31757 6307 31815 6313
rect 31757 6273 31769 6307
rect 31803 6304 31815 6307
rect 31846 6304 31852 6316
rect 31803 6276 31852 6304
rect 31803 6273 31815 6276
rect 31757 6267 31815 6273
rect 31846 6264 31852 6276
rect 31904 6264 31910 6316
rect 31956 6304 31984 6344
rect 32030 6332 32036 6384
rect 32088 6372 32094 6384
rect 33689 6375 33747 6381
rect 33689 6372 33701 6375
rect 32088 6344 33701 6372
rect 32088 6332 32094 6344
rect 33689 6341 33701 6344
rect 33735 6341 33747 6375
rect 33689 6335 33747 6341
rect 34330 6304 34336 6316
rect 31956 6276 34336 6304
rect 34330 6264 34336 6276
rect 34388 6264 34394 6316
rect 34698 6304 34704 6316
rect 34611 6276 34704 6304
rect 24578 6196 24584 6248
rect 24636 6236 24642 6248
rect 25133 6239 25191 6245
rect 25133 6236 25145 6239
rect 24636 6208 25145 6236
rect 24636 6196 24642 6208
rect 25133 6205 25145 6208
rect 25179 6205 25191 6239
rect 25133 6199 25191 6205
rect 27706 6196 27712 6248
rect 27764 6236 27770 6248
rect 27801 6239 27859 6245
rect 27801 6236 27813 6239
rect 27764 6208 27813 6236
rect 27764 6196 27770 6208
rect 27801 6205 27813 6208
rect 27847 6205 27859 6239
rect 27801 6199 27859 6205
rect 32122 6196 32128 6248
rect 32180 6236 32186 6248
rect 32180 6208 32812 6236
rect 32180 6196 32186 6208
rect 19058 6128 19064 6180
rect 19116 6168 19122 6180
rect 20165 6171 20223 6177
rect 20165 6168 20177 6171
rect 19116 6140 20177 6168
rect 19116 6128 19122 6140
rect 20165 6137 20177 6140
rect 20211 6137 20223 6171
rect 20165 6131 20223 6137
rect 22094 6128 22100 6180
rect 22152 6168 22158 6180
rect 23201 6171 23259 6177
rect 23201 6168 23213 6171
rect 22152 6140 23213 6168
rect 22152 6128 22158 6140
rect 23201 6137 23213 6140
rect 23247 6137 23259 6171
rect 23201 6131 23259 6137
rect 24946 6128 24952 6180
rect 25004 6168 25010 6180
rect 25409 6171 25467 6177
rect 25409 6168 25421 6171
rect 25004 6140 25421 6168
rect 25004 6128 25010 6140
rect 25409 6137 25421 6140
rect 25455 6137 25467 6171
rect 27430 6168 27436 6180
rect 26634 6140 27436 6168
rect 25409 6131 25467 6137
rect 27430 6128 27436 6140
rect 27488 6128 27494 6180
rect 28074 6168 28080 6180
rect 28035 6140 28080 6168
rect 28074 6128 28080 6140
rect 28132 6128 28138 6180
rect 30190 6168 30196 6180
rect 29302 6140 30196 6168
rect 30190 6128 30196 6140
rect 30248 6128 30254 6180
rect 31018 6128 31024 6180
rect 31076 6128 31082 6180
rect 31478 6168 31484 6180
rect 31439 6140 31484 6168
rect 31478 6128 31484 6140
rect 31536 6128 31542 6180
rect 32784 6168 32812 6208
rect 32950 6196 32956 6248
rect 33008 6236 33014 6248
rect 33229 6239 33287 6245
rect 33229 6236 33241 6239
rect 33008 6208 33241 6236
rect 33008 6196 33014 6208
rect 33229 6205 33241 6208
rect 33275 6205 33287 6239
rect 33870 6236 33876 6248
rect 33831 6208 33876 6236
rect 33229 6199 33287 6205
rect 33870 6196 33876 6208
rect 33928 6196 33934 6248
rect 34525 6239 34583 6245
rect 34525 6205 34537 6239
rect 34571 6236 34583 6239
rect 34624 6236 34652 6276
rect 34698 6264 34704 6276
rect 34756 6304 34762 6316
rect 35526 6304 35532 6316
rect 34756 6276 35532 6304
rect 34756 6264 34762 6276
rect 35526 6264 35532 6276
rect 35584 6264 35590 6316
rect 34571 6208 34652 6236
rect 34977 6239 35035 6245
rect 34571 6205 34583 6208
rect 34525 6199 34583 6205
rect 34977 6205 34989 6239
rect 35023 6236 35035 6239
rect 35342 6236 35348 6248
rect 35023 6208 35348 6236
rect 35023 6205 35035 6208
rect 34977 6199 35035 6205
rect 35342 6196 35348 6208
rect 35400 6196 35406 6248
rect 36078 6168 36084 6180
rect 32784 6140 36084 6168
rect 36078 6128 36084 6140
rect 36136 6128 36142 6180
rect 18690 6060 18696 6112
rect 18748 6100 18754 6112
rect 19245 6103 19303 6109
rect 19245 6100 19257 6103
rect 18748 6072 19257 6100
rect 18748 6060 18754 6072
rect 19245 6069 19257 6072
rect 19291 6069 19303 6103
rect 19245 6063 19303 6069
rect 21637 6103 21695 6109
rect 21637 6069 21649 6103
rect 21683 6100 21695 6103
rect 28810 6100 28816 6112
rect 21683 6072 28816 6100
rect 21683 6069 21695 6072
rect 21637 6063 21695 6069
rect 28810 6060 28816 6072
rect 28868 6060 28874 6112
rect 30098 6060 30104 6112
rect 30156 6100 30162 6112
rect 33045 6103 33103 6109
rect 33045 6100 33057 6103
rect 30156 6072 33057 6100
rect 30156 6060 30162 6072
rect 33045 6069 33057 6072
rect 33091 6069 33103 6103
rect 33045 6063 33103 6069
rect 35069 6103 35127 6109
rect 35069 6069 35081 6103
rect 35115 6100 35127 6103
rect 36722 6100 36728 6112
rect 35115 6072 36728 6100
rect 35115 6069 35127 6072
rect 35069 6063 35127 6069
rect 36722 6060 36728 6072
rect 36780 6060 36786 6112
rect 1104 6010 38824 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 38824 6010
rect 1104 5936 38824 5958
rect 18417 5899 18475 5905
rect 18417 5865 18429 5899
rect 18463 5896 18475 5899
rect 21358 5896 21364 5908
rect 18463 5868 21364 5896
rect 18463 5865 18475 5868
rect 18417 5859 18475 5865
rect 21358 5856 21364 5868
rect 21416 5856 21422 5908
rect 24305 5899 24363 5905
rect 21836 5868 24256 5896
rect 20070 5828 20076 5840
rect 17604 5800 20076 5828
rect 15562 5720 15568 5772
rect 15620 5760 15626 5772
rect 17604 5769 17632 5800
rect 20070 5788 20076 5800
rect 20128 5788 20134 5840
rect 21836 5814 21864 5868
rect 24118 5828 24124 5840
rect 24058 5800 24124 5828
rect 24118 5788 24124 5800
rect 24176 5788 24182 5840
rect 24228 5828 24256 5868
rect 24305 5865 24317 5899
rect 24351 5896 24363 5899
rect 24854 5896 24860 5908
rect 24351 5868 24860 5896
rect 24351 5865 24363 5868
rect 24305 5859 24363 5865
rect 24854 5856 24860 5868
rect 24912 5856 24918 5908
rect 30098 5896 30104 5908
rect 24964 5868 30104 5896
rect 24964 5828 24992 5868
rect 30098 5856 30104 5868
rect 30156 5856 30162 5908
rect 30282 5856 30288 5908
rect 30340 5896 30346 5908
rect 30469 5899 30527 5905
rect 30469 5896 30481 5899
rect 30340 5868 30481 5896
rect 30340 5856 30346 5868
rect 30469 5865 30481 5868
rect 30515 5865 30527 5899
rect 31570 5896 31576 5908
rect 30469 5859 30527 5865
rect 30668 5868 31576 5896
rect 30668 5828 30696 5868
rect 31570 5856 31576 5868
rect 31628 5856 31634 5908
rect 33042 5856 33048 5908
rect 33100 5896 33106 5908
rect 33965 5899 34023 5905
rect 33965 5896 33977 5899
rect 33100 5868 33977 5896
rect 33100 5856 33106 5868
rect 33965 5865 33977 5868
rect 34011 5865 34023 5899
rect 35710 5896 35716 5908
rect 35671 5868 35716 5896
rect 33965 5859 34023 5865
rect 35710 5856 35716 5868
rect 35768 5856 35774 5908
rect 24228 5800 24992 5828
rect 28014 5800 30696 5828
rect 31846 5788 31852 5840
rect 31904 5828 31910 5840
rect 31904 5800 32352 5828
rect 31904 5788 31910 5800
rect 17589 5763 17647 5769
rect 17589 5760 17601 5763
rect 15620 5732 17601 5760
rect 15620 5720 15626 5732
rect 17589 5729 17601 5732
rect 17635 5729 17647 5763
rect 18230 5760 18236 5772
rect 18191 5732 18236 5760
rect 17589 5723 17647 5729
rect 18230 5720 18236 5732
rect 18288 5720 18294 5772
rect 19061 5763 19119 5769
rect 19061 5729 19073 5763
rect 19107 5760 19119 5763
rect 20254 5760 20260 5772
rect 19107 5732 20260 5760
rect 19107 5729 19119 5732
rect 19061 5723 19119 5729
rect 20254 5720 20260 5732
rect 20312 5720 20318 5772
rect 22554 5760 22560 5772
rect 22515 5732 22560 5760
rect 22554 5720 22560 5732
rect 22612 5720 22618 5772
rect 25501 5763 25559 5769
rect 25501 5760 25513 5763
rect 24504 5732 25513 5760
rect 19886 5652 19892 5704
rect 19944 5692 19950 5704
rect 20349 5695 20407 5701
rect 20349 5692 20361 5695
rect 19944 5664 20361 5692
rect 19944 5652 19950 5664
rect 20349 5661 20361 5664
rect 20395 5661 20407 5695
rect 20622 5692 20628 5704
rect 20583 5664 20628 5692
rect 20349 5655 20407 5661
rect 20622 5652 20628 5664
rect 20680 5652 20686 5704
rect 22833 5695 22891 5701
rect 22833 5692 22845 5695
rect 22664 5664 22845 5692
rect 21634 5584 21640 5636
rect 21692 5624 21698 5636
rect 22664 5624 22692 5664
rect 22833 5661 22845 5664
rect 22879 5661 22891 5695
rect 22833 5655 22891 5661
rect 23382 5652 23388 5704
rect 23440 5692 23446 5704
rect 24504 5692 24532 5732
rect 25501 5729 25513 5732
rect 25547 5760 25559 5763
rect 25777 5763 25835 5769
rect 25777 5760 25789 5763
rect 25547 5732 25789 5760
rect 25547 5729 25559 5732
rect 25501 5723 25559 5729
rect 25777 5729 25789 5732
rect 25823 5729 25835 5763
rect 25777 5723 25835 5729
rect 26513 5763 26571 5769
rect 26513 5729 26525 5763
rect 26559 5760 26571 5763
rect 27154 5760 27160 5772
rect 26559 5732 27160 5760
rect 26559 5729 26571 5732
rect 26513 5723 26571 5729
rect 27154 5720 27160 5732
rect 27212 5720 27218 5772
rect 28994 5720 29000 5772
rect 29052 5760 29058 5772
rect 29181 5763 29239 5769
rect 29181 5760 29193 5763
rect 29052 5732 29193 5760
rect 29052 5720 29058 5732
rect 29181 5729 29193 5732
rect 29227 5729 29239 5763
rect 29181 5723 29239 5729
rect 30374 5720 30380 5772
rect 30432 5760 30438 5772
rect 30432 5732 30866 5760
rect 30432 5720 30438 5732
rect 25406 5692 25412 5704
rect 23440 5664 24532 5692
rect 25367 5664 25412 5692
rect 23440 5652 23446 5664
rect 25406 5652 25412 5664
rect 25464 5692 25470 5704
rect 25866 5692 25872 5704
rect 25464 5664 25872 5692
rect 25464 5652 25470 5664
rect 25866 5652 25872 5664
rect 25924 5652 25930 5704
rect 28074 5692 28080 5704
rect 25976 5664 28080 5692
rect 21692 5596 22692 5624
rect 21692 5584 21698 5596
rect 24302 5584 24308 5636
rect 24360 5624 24366 5636
rect 25976 5624 26004 5664
rect 28074 5652 28080 5664
rect 28132 5652 28138 5704
rect 28442 5692 28448 5704
rect 28403 5664 28448 5692
rect 28442 5652 28448 5664
rect 28500 5652 28506 5704
rect 28721 5695 28779 5701
rect 28721 5661 28733 5695
rect 28767 5661 28779 5695
rect 28721 5655 28779 5661
rect 24360 5596 26004 5624
rect 26329 5627 26387 5633
rect 24360 5584 24366 5596
rect 26329 5593 26341 5627
rect 26375 5624 26387 5627
rect 27430 5624 27436 5636
rect 26375 5596 27436 5624
rect 26375 5593 26387 5596
rect 26329 5587 26387 5593
rect 27430 5584 27436 5596
rect 27488 5584 27494 5636
rect 28736 5624 28764 5655
rect 28810 5652 28816 5704
rect 28868 5692 28874 5704
rect 31941 5695 31999 5701
rect 31941 5692 31953 5695
rect 28868 5664 31953 5692
rect 28868 5652 28874 5664
rect 31941 5661 31953 5664
rect 31987 5661 31999 5695
rect 32214 5692 32220 5704
rect 32175 5664 32220 5692
rect 31941 5655 31999 5661
rect 32214 5652 32220 5664
rect 32272 5652 32278 5704
rect 32324 5692 32352 5800
rect 32766 5788 32772 5840
rect 32824 5828 32830 5840
rect 33870 5828 33876 5840
rect 32824 5800 33876 5828
rect 32824 5788 32830 5800
rect 33870 5788 33876 5800
rect 33928 5828 33934 5840
rect 33928 5800 34836 5828
rect 33928 5788 33934 5800
rect 32858 5760 32864 5772
rect 32819 5732 32864 5760
rect 32858 5720 32864 5732
rect 32916 5720 32922 5772
rect 32950 5720 32956 5772
rect 33008 5760 33014 5772
rect 34808 5769 34836 5800
rect 33505 5763 33563 5769
rect 33505 5760 33517 5763
rect 33008 5732 33517 5760
rect 33008 5720 33014 5732
rect 33505 5729 33517 5732
rect 33551 5729 33563 5763
rect 33505 5723 33563 5729
rect 34149 5763 34207 5769
rect 34149 5729 34161 5763
rect 34195 5729 34207 5763
rect 34149 5723 34207 5729
rect 34793 5763 34851 5769
rect 34793 5729 34805 5763
rect 34839 5729 34851 5763
rect 35894 5760 35900 5772
rect 35855 5732 35900 5760
rect 34793 5723 34851 5729
rect 34164 5692 34192 5723
rect 32324 5664 34192 5692
rect 34808 5692 34836 5723
rect 35894 5720 35900 5732
rect 35952 5720 35958 5772
rect 36814 5692 36820 5704
rect 34808 5664 36820 5692
rect 36814 5652 36820 5664
rect 36872 5652 36878 5704
rect 30006 5624 30012 5636
rect 28736 5596 30012 5624
rect 17405 5559 17463 5565
rect 17405 5525 17417 5559
rect 17451 5556 17463 5559
rect 17494 5556 17500 5568
rect 17451 5528 17500 5556
rect 17451 5525 17463 5528
rect 17405 5519 17463 5525
rect 17494 5516 17500 5528
rect 17552 5516 17558 5568
rect 18874 5556 18880 5568
rect 18835 5528 18880 5556
rect 18874 5516 18880 5528
rect 18932 5516 18938 5568
rect 21174 5516 21180 5568
rect 21232 5556 21238 5568
rect 22097 5559 22155 5565
rect 22097 5556 22109 5559
rect 21232 5528 22109 5556
rect 21232 5516 21238 5528
rect 22097 5525 22109 5528
rect 22143 5525 22155 5559
rect 22097 5519 22155 5525
rect 24026 5516 24032 5568
rect 24084 5556 24090 5568
rect 25225 5559 25283 5565
rect 25225 5556 25237 5559
rect 24084 5528 25237 5556
rect 24084 5516 24090 5528
rect 25225 5525 25237 5528
rect 25271 5525 25283 5559
rect 25225 5519 25283 5525
rect 26973 5559 27031 5565
rect 26973 5525 26985 5559
rect 27019 5556 27031 5559
rect 27798 5556 27804 5568
rect 27019 5528 27804 5556
rect 27019 5525 27031 5528
rect 26973 5519 27031 5525
rect 27798 5516 27804 5528
rect 27856 5516 27862 5568
rect 27982 5516 27988 5568
rect 28040 5556 28046 5568
rect 28736 5556 28764 5596
rect 30006 5584 30012 5596
rect 30064 5584 30070 5636
rect 30190 5584 30196 5636
rect 30248 5624 30254 5636
rect 34609 5627 34667 5633
rect 34609 5624 34621 5627
rect 30248 5596 30604 5624
rect 30248 5584 30254 5596
rect 29362 5556 29368 5568
rect 28040 5528 28764 5556
rect 29323 5528 29368 5556
rect 28040 5516 28046 5528
rect 29362 5516 29368 5528
rect 29420 5556 29426 5568
rect 29822 5556 29828 5568
rect 29420 5528 29828 5556
rect 29420 5516 29426 5528
rect 29822 5516 29828 5528
rect 29880 5516 29886 5568
rect 30576 5556 30604 5596
rect 32600 5596 34621 5624
rect 32600 5556 32628 5596
rect 34609 5593 34621 5596
rect 34655 5593 34667 5627
rect 34609 5587 34667 5593
rect 30576 5528 32628 5556
rect 32677 5559 32735 5565
rect 32677 5525 32689 5559
rect 32723 5556 32735 5559
rect 32766 5556 32772 5568
rect 32723 5528 32772 5556
rect 32723 5525 32735 5528
rect 32677 5519 32735 5525
rect 32766 5516 32772 5528
rect 32824 5516 32830 5568
rect 33318 5556 33324 5568
rect 33279 5528 33324 5556
rect 33318 5516 33324 5528
rect 33376 5516 33382 5568
rect 33410 5516 33416 5568
rect 33468 5556 33474 5568
rect 36446 5556 36452 5568
rect 33468 5528 36452 5556
rect 33468 5516 33474 5528
rect 36446 5516 36452 5528
rect 36504 5516 36510 5568
rect 1104 5466 38824 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 38824 5466
rect 1104 5392 38824 5414
rect 17310 5312 17316 5364
rect 17368 5352 17374 5364
rect 19165 5355 19223 5361
rect 19165 5352 19177 5355
rect 17368 5324 19177 5352
rect 17368 5312 17374 5324
rect 19165 5321 19177 5324
rect 19211 5352 19223 5355
rect 19334 5352 19340 5364
rect 19211 5324 19340 5352
rect 19211 5321 19223 5324
rect 19165 5315 19223 5321
rect 19334 5312 19340 5324
rect 19392 5312 19398 5364
rect 21637 5355 21695 5361
rect 21637 5321 21649 5355
rect 21683 5352 21695 5355
rect 21726 5352 21732 5364
rect 21683 5324 21732 5352
rect 21683 5321 21695 5324
rect 21637 5315 21695 5321
rect 21726 5312 21732 5324
rect 21784 5312 21790 5364
rect 23106 5312 23112 5364
rect 23164 5352 23170 5364
rect 31757 5355 31815 5361
rect 31757 5352 31769 5355
rect 23164 5324 31769 5352
rect 23164 5312 23170 5324
rect 31757 5321 31769 5324
rect 31803 5321 31815 5355
rect 31757 5315 31815 5321
rect 35710 5312 35716 5364
rect 35768 5352 35774 5364
rect 35897 5355 35955 5361
rect 35897 5352 35909 5355
rect 35768 5324 35909 5352
rect 35768 5312 35774 5324
rect 35897 5321 35909 5324
rect 35943 5321 35955 5355
rect 35897 5315 35955 5321
rect 25130 5284 25136 5296
rect 24688 5256 25136 5284
rect 17494 5176 17500 5228
rect 17552 5216 17558 5228
rect 19429 5219 19487 5225
rect 19429 5216 19441 5219
rect 17552 5188 19441 5216
rect 17552 5176 17558 5188
rect 19429 5185 19441 5188
rect 19475 5216 19487 5219
rect 19886 5216 19892 5228
rect 19475 5188 19892 5216
rect 19475 5185 19487 5188
rect 19429 5179 19487 5185
rect 19886 5176 19892 5188
rect 19944 5176 19950 5228
rect 20165 5219 20223 5225
rect 20165 5185 20177 5219
rect 20211 5216 20223 5219
rect 21174 5216 21180 5228
rect 20211 5188 21180 5216
rect 20211 5185 20223 5188
rect 20165 5179 20223 5185
rect 21174 5176 21180 5188
rect 21232 5176 21238 5228
rect 22830 5216 22836 5228
rect 21284 5188 22836 5216
rect 21284 5134 21312 5188
rect 22830 5176 22836 5188
rect 22888 5176 22894 5228
rect 24688 5225 24716 5256
rect 25130 5244 25136 5256
rect 25188 5244 25194 5296
rect 29638 5284 29644 5296
rect 29472 5256 29644 5284
rect 24673 5219 24731 5225
rect 24673 5216 24685 5219
rect 23216 5188 24685 5216
rect 22462 5108 22468 5160
rect 22520 5148 22526 5160
rect 23216 5148 23244 5188
rect 24673 5185 24685 5188
rect 24719 5185 24731 5219
rect 24673 5179 24731 5185
rect 27430 5176 27436 5228
rect 27488 5216 27494 5228
rect 28810 5216 28816 5228
rect 27488 5188 28816 5216
rect 27488 5176 27494 5188
rect 28810 5176 28816 5188
rect 28868 5176 28874 5228
rect 29273 5219 29331 5225
rect 29273 5185 29285 5219
rect 29319 5216 29331 5219
rect 29472 5216 29500 5256
rect 29638 5244 29644 5256
rect 29696 5244 29702 5296
rect 33042 5284 33048 5296
rect 31312 5256 33048 5284
rect 29319 5188 29500 5216
rect 29319 5185 29331 5188
rect 29273 5179 29331 5185
rect 29546 5176 29552 5228
rect 29604 5216 29610 5228
rect 29604 5188 29649 5216
rect 29604 5176 29610 5188
rect 29730 5176 29736 5228
rect 29788 5216 29794 5228
rect 31312 5216 31340 5256
rect 33042 5244 33048 5256
rect 33100 5244 33106 5296
rect 34793 5287 34851 5293
rect 34793 5253 34805 5287
rect 34839 5284 34851 5287
rect 35986 5284 35992 5296
rect 34839 5256 35992 5284
rect 34839 5253 34851 5256
rect 34793 5247 34851 5253
rect 35986 5244 35992 5256
rect 36044 5244 36050 5296
rect 36541 5287 36599 5293
rect 36541 5253 36553 5287
rect 36587 5253 36599 5287
rect 36541 5247 36599 5253
rect 36556 5216 36584 5247
rect 29788 5188 31340 5216
rect 32140 5188 36584 5216
rect 29788 5176 29794 5188
rect 25130 5148 25136 5160
rect 22520 5120 23244 5148
rect 25091 5120 25136 5148
rect 22520 5108 22526 5120
rect 25130 5108 25136 5120
rect 25188 5108 25194 5160
rect 29564 5148 29592 5176
rect 30009 5151 30067 5157
rect 30009 5148 30021 5151
rect 29564 5120 30021 5148
rect 30009 5117 30021 5120
rect 30055 5117 30067 5151
rect 30009 5111 30067 5117
rect 20438 5080 20444 5092
rect 18722 5052 20444 5080
rect 20438 5040 20444 5052
rect 20496 5040 20502 5092
rect 22830 5080 22836 5092
rect 21468 5052 22836 5080
rect 15194 4972 15200 5024
rect 15252 5012 15258 5024
rect 17681 5015 17739 5021
rect 17681 5012 17693 5015
rect 15252 4984 17693 5012
rect 15252 4972 15258 4984
rect 17681 4981 17693 4984
rect 17727 4981 17739 5015
rect 17681 4975 17739 4981
rect 19978 4972 19984 5024
rect 20036 5012 20042 5024
rect 21468 5012 21496 5052
rect 22830 5040 22836 5052
rect 22888 5040 22894 5092
rect 23658 5040 23664 5092
rect 23716 5040 23722 5092
rect 24118 5040 24124 5092
rect 24176 5080 24182 5092
rect 24397 5083 24455 5089
rect 24397 5080 24409 5083
rect 24176 5052 24409 5080
rect 24176 5040 24182 5052
rect 24397 5049 24409 5052
rect 24443 5049 24455 5083
rect 25406 5080 25412 5092
rect 25367 5052 25412 5080
rect 24397 5043 24455 5049
rect 25406 5040 25412 5052
rect 25464 5040 25470 5092
rect 27522 5080 27528 5092
rect 26634 5052 27528 5080
rect 27522 5040 27528 5052
rect 27580 5040 27586 5092
rect 20036 4984 21496 5012
rect 20036 4972 20042 4984
rect 21542 4972 21548 5024
rect 21600 5012 21606 5024
rect 22925 5015 22983 5021
rect 22925 5012 22937 5015
rect 21600 4984 22937 5012
rect 21600 4972 21606 4984
rect 22925 4981 22937 4984
rect 22971 4981 22983 5015
rect 22925 4975 22983 4981
rect 25498 4972 25504 5024
rect 25556 5012 25562 5024
rect 26881 5015 26939 5021
rect 26881 5012 26893 5015
rect 25556 4984 26893 5012
rect 25556 4972 25562 4984
rect 26881 4981 26893 4984
rect 26927 4981 26939 5015
rect 26881 4975 26939 4981
rect 27706 4972 27712 5024
rect 27764 5012 27770 5024
rect 27801 5015 27859 5021
rect 27801 5012 27813 5015
rect 27764 4984 27813 5012
rect 27764 4972 27770 4984
rect 27801 4981 27813 4984
rect 27847 4981 27859 5015
rect 28828 5012 28856 5066
rect 28994 5040 29000 5092
rect 29052 5080 29058 5092
rect 30285 5083 30343 5089
rect 30285 5080 30297 5083
rect 29052 5052 30297 5080
rect 29052 5040 29058 5052
rect 30285 5049 30297 5052
rect 30331 5049 30343 5083
rect 30285 5043 30343 5049
rect 30374 5040 30380 5092
rect 30432 5080 30438 5092
rect 30558 5080 30564 5092
rect 30432 5052 30564 5080
rect 30432 5040 30438 5052
rect 30558 5040 30564 5052
rect 30616 5040 30622 5092
rect 31294 5040 31300 5092
rect 31352 5040 31358 5092
rect 32140 5012 32168 5188
rect 32214 5108 32220 5160
rect 32272 5148 32278 5160
rect 33042 5148 33048 5160
rect 32272 5120 33048 5148
rect 32272 5108 32278 5120
rect 33042 5108 33048 5120
rect 33100 5108 33106 5160
rect 35434 5148 35440 5160
rect 35395 5120 35440 5148
rect 35434 5108 35440 5120
rect 35492 5108 35498 5160
rect 35526 5108 35532 5160
rect 35584 5148 35590 5160
rect 36081 5151 36139 5157
rect 36081 5148 36093 5151
rect 35584 5120 36093 5148
rect 35584 5108 35590 5120
rect 36081 5117 36093 5120
rect 36127 5117 36139 5151
rect 36081 5111 36139 5117
rect 36725 5151 36783 5157
rect 36725 5117 36737 5151
rect 36771 5117 36783 5151
rect 36725 5111 36783 5117
rect 32490 5040 32496 5092
rect 32548 5080 32554 5092
rect 33321 5083 33379 5089
rect 33321 5080 33333 5083
rect 32548 5052 33333 5080
rect 32548 5040 32554 5052
rect 33321 5049 33333 5052
rect 33367 5049 33379 5083
rect 33321 5043 33379 5049
rect 33778 5040 33784 5092
rect 33836 5040 33842 5092
rect 35894 5040 35900 5092
rect 35952 5080 35958 5092
rect 36740 5080 36768 5111
rect 35952 5052 36768 5080
rect 35952 5040 35958 5052
rect 28828 4984 32168 5012
rect 27801 4975 27859 4981
rect 32214 4972 32220 5024
rect 32272 5012 32278 5024
rect 34238 5012 34244 5024
rect 32272 4984 34244 5012
rect 32272 4972 32278 4984
rect 34238 4972 34244 4984
rect 34296 4972 34302 5024
rect 34330 4972 34336 5024
rect 34388 5012 34394 5024
rect 35253 5015 35311 5021
rect 35253 5012 35265 5015
rect 34388 4984 35265 5012
rect 34388 4972 34394 4984
rect 35253 4981 35265 4984
rect 35299 4981 35311 5015
rect 35253 4975 35311 4981
rect 1104 4922 38824 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 38824 4922
rect 1104 4848 38824 4870
rect 18874 4808 18880 4820
rect 16684 4780 18880 4808
rect 16684 4681 16712 4780
rect 18874 4768 18880 4780
rect 18932 4768 18938 4820
rect 19334 4768 19340 4820
rect 19392 4808 19398 4820
rect 21450 4808 21456 4820
rect 19392 4780 21456 4808
rect 19392 4768 19398 4780
rect 21450 4768 21456 4780
rect 21508 4768 21514 4820
rect 35713 4811 35771 4817
rect 35713 4808 35725 4811
rect 21836 4780 35725 4808
rect 17494 4740 17500 4752
rect 17328 4712 17500 4740
rect 17328 4681 17356 4712
rect 17494 4700 17500 4712
rect 17552 4700 17558 4752
rect 21836 4726 21864 4780
rect 35713 4777 35725 4780
rect 35759 4777 35771 4811
rect 35713 4771 35771 4777
rect 35802 4768 35808 4820
rect 35860 4808 35866 4820
rect 37645 4811 37703 4817
rect 37645 4808 37657 4811
rect 35860 4780 37657 4808
rect 35860 4768 35866 4780
rect 37645 4777 37657 4780
rect 37691 4777 37703 4811
rect 37645 4771 37703 4777
rect 23106 4740 23112 4752
rect 21928 4712 23112 4740
rect 16669 4675 16727 4681
rect 16669 4641 16681 4675
rect 16715 4641 16727 4675
rect 16669 4635 16727 4641
rect 17313 4675 17371 4681
rect 17313 4641 17325 4675
rect 17359 4641 17371 4675
rect 18722 4644 20116 4672
rect 17313 4635 17371 4641
rect 17586 4604 17592 4616
rect 17547 4576 17592 4604
rect 17586 4564 17592 4576
rect 17644 4564 17650 4616
rect 16853 4471 16911 4477
rect 16853 4437 16865 4471
rect 16899 4468 16911 4471
rect 18046 4468 18052 4480
rect 16899 4440 18052 4468
rect 16899 4437 16911 4440
rect 16853 4431 16911 4437
rect 18046 4428 18052 4440
rect 18104 4428 18110 4480
rect 19061 4471 19119 4477
rect 19061 4437 19073 4471
rect 19107 4468 19119 4471
rect 19150 4468 19156 4480
rect 19107 4440 19156 4468
rect 19107 4437 19119 4440
rect 19061 4431 19119 4437
rect 19150 4428 19156 4440
rect 19208 4428 19214 4480
rect 20088 4468 20116 4644
rect 20346 4604 20352 4616
rect 20307 4576 20352 4604
rect 20346 4564 20352 4576
rect 20404 4564 20410 4616
rect 20625 4607 20683 4613
rect 20625 4573 20637 4607
rect 20671 4604 20683 4607
rect 21928 4604 21956 4712
rect 23106 4700 23112 4712
rect 23164 4700 23170 4752
rect 25498 4740 25504 4752
rect 25459 4712 25504 4740
rect 25498 4700 25504 4712
rect 25556 4700 25562 4752
rect 27430 4740 27436 4752
rect 26726 4712 27436 4740
rect 27430 4700 27436 4712
rect 27488 4700 27494 4752
rect 27706 4740 27712 4752
rect 27667 4712 27712 4740
rect 27706 4700 27712 4712
rect 27764 4700 27770 4752
rect 28350 4700 28356 4752
rect 28408 4700 28414 4752
rect 30006 4700 30012 4752
rect 30064 4740 30070 4752
rect 30742 4740 30748 4752
rect 30064 4712 30512 4740
rect 30703 4712 30748 4740
rect 30064 4700 30070 4712
rect 20671 4576 21956 4604
rect 20671 4573 20683 4576
rect 20625 4567 20683 4573
rect 22094 4564 22100 4616
rect 22152 4604 22158 4616
rect 22554 4604 22560 4616
rect 22152 4576 22197 4604
rect 22515 4576 22560 4604
rect 22152 4564 22158 4576
rect 22554 4564 22560 4576
rect 22612 4564 22618 4616
rect 22830 4604 22836 4616
rect 22791 4576 22836 4604
rect 22830 4564 22836 4576
rect 22888 4564 22894 4616
rect 23198 4564 23204 4616
rect 23256 4604 23262 4616
rect 23474 4604 23480 4616
rect 23256 4576 23480 4604
rect 23256 4564 23262 4576
rect 23474 4564 23480 4576
rect 23532 4564 23538 4616
rect 23952 4604 23980 4658
rect 25130 4632 25136 4684
rect 25188 4672 25194 4684
rect 25225 4675 25283 4681
rect 25225 4672 25237 4675
rect 25188 4644 25237 4672
rect 25188 4632 25194 4644
rect 25225 4641 25237 4644
rect 25271 4641 25283 4675
rect 30374 4672 30380 4684
rect 25225 4635 25283 4641
rect 28920 4644 30380 4672
rect 27430 4604 27436 4616
rect 23952 4576 26556 4604
rect 27391 4576 27436 4604
rect 26528 4536 26556 4576
rect 27430 4564 27436 4576
rect 27488 4564 27494 4616
rect 28920 4604 28948 4644
rect 30374 4632 30380 4644
rect 30432 4632 30438 4684
rect 30484 4681 30512 4712
rect 30742 4700 30748 4712
rect 30800 4700 30806 4752
rect 32858 4740 32864 4752
rect 31970 4712 32864 4740
rect 32858 4700 32864 4712
rect 32916 4700 32922 4752
rect 35250 4740 35256 4752
rect 33718 4712 35256 4740
rect 35250 4700 35256 4712
rect 35308 4700 35314 4752
rect 30469 4675 30527 4681
rect 30469 4641 30481 4675
rect 30515 4641 30527 4675
rect 30469 4635 30527 4641
rect 34514 4632 34520 4684
rect 34572 4672 34578 4684
rect 35342 4672 35348 4684
rect 34572 4644 35348 4672
rect 34572 4632 34578 4644
rect 35342 4632 35348 4644
rect 35400 4632 35406 4684
rect 35434 4632 35440 4684
rect 35492 4672 35498 4684
rect 35897 4675 35955 4681
rect 35897 4672 35909 4675
rect 35492 4644 35909 4672
rect 35492 4632 35498 4644
rect 35897 4641 35909 4644
rect 35943 4672 35955 4675
rect 36354 4672 36360 4684
rect 35943 4644 36360 4672
rect 35943 4641 35955 4644
rect 35897 4635 35955 4641
rect 36354 4632 36360 4644
rect 36412 4632 36418 4684
rect 36541 4675 36599 4681
rect 36541 4641 36553 4675
rect 36587 4672 36599 4675
rect 36814 4672 36820 4684
rect 36587 4644 36820 4672
rect 36587 4641 36599 4644
rect 36541 4635 36599 4641
rect 36814 4632 36820 4644
rect 36872 4632 36878 4684
rect 37185 4675 37243 4681
rect 37185 4641 37197 4675
rect 37231 4641 37243 4675
rect 37826 4672 37832 4684
rect 37787 4644 37832 4672
rect 37185 4635 37243 4641
rect 29178 4604 29184 4616
rect 27540 4576 28948 4604
rect 29139 4576 29184 4604
rect 27540 4536 27568 4576
rect 29178 4564 29184 4576
rect 29236 4564 29242 4616
rect 31478 4604 31484 4616
rect 30208 4576 31484 4604
rect 30208 4536 30236 4576
rect 31478 4564 31484 4576
rect 31536 4564 31542 4616
rect 34146 4604 34152 4616
rect 34107 4576 34152 4604
rect 34146 4564 34152 4576
rect 34204 4564 34210 4616
rect 34425 4607 34483 4613
rect 34425 4573 34437 4607
rect 34471 4604 34483 4607
rect 34606 4604 34612 4616
rect 34471 4576 34612 4604
rect 34471 4573 34483 4576
rect 34425 4567 34483 4573
rect 34606 4564 34612 4576
rect 34664 4564 34670 4616
rect 34698 4564 34704 4616
rect 34756 4604 34762 4616
rect 37200 4604 37228 4635
rect 37826 4632 37832 4644
rect 37884 4632 37890 4684
rect 34756 4576 37228 4604
rect 34756 4564 34762 4576
rect 37001 4539 37059 4545
rect 37001 4536 37013 4539
rect 26528 4508 27568 4536
rect 28736 4508 30236 4536
rect 32094 4508 32812 4536
rect 23198 4468 23204 4480
rect 20088 4440 23204 4468
rect 23198 4428 23204 4440
rect 23256 4428 23262 4480
rect 23474 4428 23480 4480
rect 23532 4468 23538 4480
rect 24305 4471 24363 4477
rect 24305 4468 24317 4471
rect 23532 4440 24317 4468
rect 23532 4428 23538 4440
rect 24305 4437 24317 4440
rect 24351 4437 24363 4471
rect 24305 4431 24363 4437
rect 26973 4471 27031 4477
rect 26973 4437 26985 4471
rect 27019 4468 27031 4471
rect 27154 4468 27160 4480
rect 27019 4440 27160 4468
rect 27019 4437 27031 4440
rect 26973 4431 27031 4437
rect 27154 4428 27160 4440
rect 27212 4428 27218 4480
rect 27706 4428 27712 4480
rect 27764 4468 27770 4480
rect 28736 4468 28764 4508
rect 27764 4440 28764 4468
rect 27764 4428 27770 4440
rect 29638 4428 29644 4480
rect 29696 4468 29702 4480
rect 32094 4468 32122 4508
rect 32214 4468 32220 4480
rect 29696 4440 32122 4468
rect 32175 4440 32220 4468
rect 29696 4428 29702 4440
rect 32214 4428 32220 4440
rect 32272 4428 32278 4480
rect 32674 4468 32680 4480
rect 32635 4440 32680 4468
rect 32674 4428 32680 4440
rect 32732 4428 32738 4480
rect 32784 4468 32812 4508
rect 34348 4508 37013 4536
rect 34348 4468 34376 4508
rect 37001 4505 37013 4508
rect 37047 4505 37059 4539
rect 37001 4499 37059 4505
rect 32784 4440 34376 4468
rect 34422 4428 34428 4480
rect 34480 4468 34486 4480
rect 36357 4471 36415 4477
rect 36357 4468 36369 4471
rect 34480 4440 36369 4468
rect 34480 4428 34486 4440
rect 36357 4437 36369 4440
rect 36403 4437 36415 4471
rect 36357 4431 36415 4437
rect 1104 4378 38824 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 38824 4378
rect 1104 4304 38824 4326
rect 17944 4267 18002 4273
rect 17944 4233 17956 4267
rect 17990 4264 18002 4267
rect 19978 4264 19984 4276
rect 17990 4236 19984 4264
rect 17990 4233 18002 4236
rect 17944 4227 18002 4233
rect 19978 4224 19984 4236
rect 20036 4224 20042 4276
rect 20152 4267 20210 4273
rect 20152 4233 20164 4267
rect 20198 4264 20210 4267
rect 23188 4267 23246 4273
rect 20198 4236 23060 4264
rect 20198 4233 20210 4236
rect 20152 4227 20210 4233
rect 21450 4156 21456 4208
rect 21508 4196 21514 4208
rect 21726 4196 21732 4208
rect 21508 4168 21732 4196
rect 21508 4156 21514 4168
rect 21726 4156 21732 4168
rect 21784 4156 21790 4208
rect 19429 4131 19487 4137
rect 19429 4097 19441 4131
rect 19475 4128 19487 4131
rect 20622 4128 20628 4140
rect 19475 4100 20628 4128
rect 19475 4097 19487 4100
rect 19429 4091 19487 4097
rect 20622 4088 20628 4100
rect 20680 4088 20686 4140
rect 21634 4128 21640 4140
rect 21595 4100 21640 4128
rect 21634 4088 21640 4100
rect 21692 4088 21698 4140
rect 22462 4088 22468 4140
rect 22520 4128 22526 4140
rect 22925 4131 22983 4137
rect 22925 4128 22937 4131
rect 22520 4100 22937 4128
rect 22520 4088 22526 4100
rect 22925 4097 22937 4100
rect 22971 4097 22983 4131
rect 23032 4128 23060 4236
rect 23188 4233 23200 4267
rect 23234 4264 23246 4267
rect 24854 4264 24860 4276
rect 23234 4236 24860 4264
rect 23234 4233 23246 4236
rect 23188 4227 23246 4233
rect 24854 4224 24860 4236
rect 24912 4224 24918 4276
rect 25133 4267 25191 4273
rect 25133 4233 25145 4267
rect 25179 4264 25191 4267
rect 25406 4264 25412 4276
rect 25179 4236 25412 4264
rect 25179 4233 25191 4236
rect 25133 4227 25191 4233
rect 25406 4224 25412 4236
rect 25464 4224 25470 4276
rect 26970 4264 26976 4276
rect 25516 4236 26976 4264
rect 25516 4196 25544 4236
rect 26970 4224 26976 4236
rect 27028 4224 27034 4276
rect 27798 4224 27804 4276
rect 27856 4264 27862 4276
rect 28058 4267 28116 4273
rect 28058 4264 28070 4267
rect 27856 4236 28070 4264
rect 27856 4224 27862 4236
rect 28058 4233 28070 4236
rect 28104 4233 28116 4267
rect 28058 4227 28116 4233
rect 28442 4224 28448 4276
rect 28500 4264 28506 4276
rect 28626 4264 28632 4276
rect 28500 4236 28632 4264
rect 28500 4224 28506 4236
rect 28626 4224 28632 4236
rect 28684 4224 28690 4276
rect 29546 4264 29552 4276
rect 29507 4236 29552 4264
rect 29546 4224 29552 4236
rect 29604 4224 29610 4276
rect 30466 4224 30472 4276
rect 30524 4264 30530 4276
rect 30524 4236 31754 4264
rect 30524 4224 30530 4236
rect 31726 4196 31754 4236
rect 33042 4224 33048 4276
rect 33100 4264 33106 4276
rect 34146 4264 34152 4276
rect 33100 4236 34152 4264
rect 33100 4224 33106 4236
rect 34146 4224 34152 4236
rect 34204 4224 34210 4276
rect 34330 4224 34336 4276
rect 34388 4264 34394 4276
rect 34698 4264 34704 4276
rect 34388 4236 34704 4264
rect 34388 4224 34394 4236
rect 34698 4224 34704 4236
rect 34756 4224 34762 4276
rect 35250 4264 35256 4276
rect 35211 4236 35256 4264
rect 35250 4224 35256 4236
rect 35308 4224 35314 4276
rect 33502 4196 33508 4208
rect 24228 4168 25544 4196
rect 26804 4168 27936 4196
rect 31726 4168 33508 4196
rect 24228 4128 24256 4168
rect 23032 4100 24256 4128
rect 26605 4131 26663 4137
rect 22925 4091 22983 4097
rect 26605 4097 26617 4131
rect 26651 4128 26663 4131
rect 26804 4128 26832 4168
rect 26651 4100 26832 4128
rect 26651 4097 26663 4100
rect 26605 4091 26663 4097
rect 26878 4088 26884 4140
rect 26936 4128 26942 4140
rect 27614 4128 27620 4140
rect 26936 4100 27620 4128
rect 26936 4088 26942 4100
rect 27614 4088 27620 4100
rect 27672 4128 27678 4140
rect 27798 4128 27804 4140
rect 27672 4100 27804 4128
rect 27672 4088 27678 4100
rect 27798 4088 27804 4100
rect 27856 4088 27862 4140
rect 27908 4128 27936 4168
rect 33502 4156 33508 4168
rect 33560 4156 33566 4208
rect 30009 4131 30067 4137
rect 30009 4128 30021 4131
rect 27908 4100 30021 4128
rect 30009 4097 30021 4100
rect 30055 4097 30067 4131
rect 30009 4091 30067 4097
rect 31478 4088 31484 4140
rect 31536 4128 31542 4140
rect 31536 4100 31581 4128
rect 31536 4088 31542 4100
rect 32030 4088 32036 4140
rect 32088 4128 32094 4140
rect 32088 4100 35480 4128
rect 32088 4088 32094 4100
rect 15562 4060 15568 4072
rect 15523 4032 15568 4060
rect 15562 4020 15568 4032
rect 15620 4020 15626 4072
rect 16209 4063 16267 4069
rect 16209 4029 16221 4063
rect 16255 4060 16267 4063
rect 17218 4060 17224 4072
rect 16255 4032 17224 4060
rect 16255 4029 16267 4032
rect 16209 4023 16267 4029
rect 17218 4020 17224 4032
rect 17276 4020 17282 4072
rect 17494 4020 17500 4072
rect 17552 4060 17558 4072
rect 17681 4063 17739 4069
rect 17681 4060 17693 4063
rect 17552 4032 17693 4060
rect 17552 4020 17558 4032
rect 17681 4029 17693 4032
rect 17727 4029 17739 4063
rect 19886 4060 19892 4072
rect 19847 4032 19892 4060
rect 17681 4023 17739 4029
rect 19886 4020 19892 4032
rect 19944 4020 19950 4072
rect 31757 4063 31815 4069
rect 31757 4029 31769 4063
rect 31803 4060 31815 4063
rect 31846 4060 31852 4072
rect 31803 4032 31852 4060
rect 31803 4029 31815 4032
rect 31757 4023 31815 4029
rect 31846 4020 31852 4032
rect 31904 4020 31910 4072
rect 34790 4020 34796 4072
rect 34848 4060 34854 4072
rect 35452 4069 35480 4100
rect 35437 4063 35495 4069
rect 34848 4032 34893 4060
rect 34848 4020 34854 4032
rect 35437 4029 35449 4063
rect 35483 4029 35495 4063
rect 36078 4060 36084 4072
rect 36039 4032 36084 4060
rect 35437 4023 35495 4029
rect 36078 4020 36084 4032
rect 36136 4020 36142 4072
rect 36354 4020 36360 4072
rect 36412 4060 36418 4072
rect 36725 4063 36783 4069
rect 36725 4060 36737 4063
rect 36412 4032 36737 4060
rect 36412 4020 36418 4032
rect 36725 4029 36737 4032
rect 36771 4029 36783 4063
rect 36725 4023 36783 4029
rect 17954 3992 17960 4004
rect 15764 3964 17960 3992
rect 15764 3933 15792 3964
rect 17954 3952 17960 3964
rect 18012 3952 18018 4004
rect 19242 3992 19248 4004
rect 19182 3964 19248 3992
rect 19242 3952 19248 3964
rect 19300 3952 19306 4004
rect 21450 3992 21456 4004
rect 21390 3964 21456 3992
rect 21450 3952 21456 3964
rect 21508 3952 21514 4004
rect 25314 3992 25320 4004
rect 24426 3964 25320 3992
rect 25314 3952 25320 3964
rect 25372 3952 25378 4004
rect 15749 3927 15807 3933
rect 15749 3893 15761 3927
rect 15795 3893 15807 3927
rect 16390 3924 16396 3936
rect 16351 3896 16396 3924
rect 15749 3887 15807 3893
rect 16390 3884 16396 3896
rect 16448 3884 16454 3936
rect 18598 3884 18604 3936
rect 18656 3924 18662 3936
rect 22186 3924 22192 3936
rect 18656 3896 22192 3924
rect 18656 3884 18662 3896
rect 22186 3884 22192 3896
rect 22244 3884 22250 3936
rect 24673 3927 24731 3933
rect 24673 3893 24685 3927
rect 24719 3924 24731 3927
rect 25682 3924 25688 3936
rect 24719 3896 25688 3924
rect 24719 3893 24731 3896
rect 24673 3887 24731 3893
rect 25682 3884 25688 3896
rect 25740 3884 25746 3936
rect 26160 3924 26188 3978
rect 28718 3952 28724 4004
rect 28776 3952 28782 4004
rect 31018 3952 31024 4004
rect 31076 3952 31082 4004
rect 31202 3952 31208 4004
rect 31260 3992 31266 4004
rect 34517 3995 34575 4001
rect 31260 3964 33350 3992
rect 31260 3952 31266 3964
rect 34517 3961 34529 3995
rect 34563 3961 34575 3995
rect 36740 3992 36768 4023
rect 36814 4020 36820 4072
rect 36872 4060 36878 4072
rect 37369 4063 37427 4069
rect 37369 4060 37381 4063
rect 36872 4032 37381 4060
rect 36872 4020 36878 4032
rect 37369 4029 37381 4032
rect 37415 4060 37427 4063
rect 37826 4060 37832 4072
rect 37415 4032 37832 4060
rect 37415 4029 37427 4032
rect 37369 4023 37427 4029
rect 37826 4020 37832 4032
rect 37884 4020 37890 4072
rect 36998 3992 37004 4004
rect 36740 3964 37004 3992
rect 34517 3955 34575 3961
rect 31570 3924 31576 3936
rect 26160 3896 31576 3924
rect 31570 3884 31576 3896
rect 31628 3884 31634 3936
rect 32398 3884 32404 3936
rect 32456 3924 32462 3936
rect 33045 3927 33103 3933
rect 33045 3924 33057 3927
rect 32456 3896 33057 3924
rect 32456 3884 32462 3896
rect 33045 3893 33057 3896
rect 33091 3893 33103 3927
rect 33045 3887 33103 3893
rect 33502 3884 33508 3936
rect 33560 3924 33566 3936
rect 34532 3924 34560 3955
rect 36998 3952 37004 3964
rect 37056 3952 37062 4004
rect 33560 3896 34560 3924
rect 33560 3884 33566 3896
rect 34606 3884 34612 3936
rect 34664 3924 34670 3936
rect 35897 3927 35955 3933
rect 35897 3924 35909 3927
rect 34664 3896 35909 3924
rect 34664 3884 34670 3896
rect 35897 3893 35909 3896
rect 35943 3893 35955 3927
rect 36538 3924 36544 3936
rect 36499 3896 36544 3924
rect 35897 3887 35955 3893
rect 36538 3884 36544 3896
rect 36596 3884 36602 3936
rect 36814 3884 36820 3936
rect 36872 3924 36878 3936
rect 37185 3927 37243 3933
rect 37185 3924 37197 3927
rect 36872 3896 37197 3924
rect 36872 3884 36878 3896
rect 37185 3893 37197 3896
rect 37231 3893 37243 3927
rect 37185 3887 37243 3893
rect 1104 3834 38824 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 38824 3834
rect 1104 3760 38824 3782
rect 18598 3720 18604 3732
rect 15396 3692 18604 3720
rect 15396 3661 15424 3692
rect 18598 3680 18604 3692
rect 18656 3680 18662 3732
rect 19058 3720 19064 3732
rect 19019 3692 19064 3720
rect 19058 3680 19064 3692
rect 19116 3680 19122 3732
rect 25225 3723 25283 3729
rect 25225 3720 25237 3723
rect 20640 3692 25237 3720
rect 15381 3655 15439 3661
rect 15381 3621 15393 3655
rect 15427 3621 15439 3655
rect 15381 3615 15439 3621
rect 16114 3612 16120 3664
rect 16172 3612 16178 3664
rect 17494 3652 17500 3664
rect 17328 3624 17500 3652
rect 14642 3476 14648 3528
rect 14700 3516 14706 3528
rect 17328 3525 17356 3624
rect 17494 3612 17500 3624
rect 17552 3612 17558 3664
rect 18046 3612 18052 3664
rect 18104 3612 18110 3664
rect 20640 3661 20668 3692
rect 25225 3689 25237 3692
rect 25271 3689 25283 3723
rect 25225 3683 25283 3689
rect 25314 3680 25320 3732
rect 25372 3720 25378 3732
rect 28442 3720 28448 3732
rect 25372 3692 28448 3720
rect 25372 3680 25378 3692
rect 28442 3680 28448 3692
rect 28500 3680 28506 3732
rect 28626 3720 28632 3732
rect 28587 3692 28632 3720
rect 28626 3680 28632 3692
rect 28684 3680 28690 3732
rect 28718 3680 28724 3732
rect 28776 3720 28782 3732
rect 31202 3720 31208 3732
rect 28776 3692 31208 3720
rect 28776 3680 28782 3692
rect 31202 3680 31208 3692
rect 31260 3680 31266 3732
rect 36814 3720 36820 3732
rect 31772 3692 36820 3720
rect 20625 3655 20683 3661
rect 20625 3621 20637 3655
rect 20671 3621 20683 3655
rect 21910 3652 21916 3664
rect 21850 3624 21916 3652
rect 20625 3615 20683 3621
rect 21910 3612 21916 3624
rect 21968 3612 21974 3664
rect 22833 3655 22891 3661
rect 22833 3621 22845 3655
rect 22879 3652 22891 3655
rect 22922 3652 22928 3664
rect 22879 3624 22928 3652
rect 22879 3621 22891 3624
rect 22833 3615 22891 3621
rect 22922 3612 22928 3624
rect 22980 3612 22986 3664
rect 25774 3652 25780 3664
rect 25516 3624 25780 3652
rect 22554 3584 22560 3596
rect 21836 3556 22560 3584
rect 15105 3519 15163 3525
rect 15105 3516 15117 3519
rect 14700 3488 15117 3516
rect 14700 3476 14706 3488
rect 15105 3485 15117 3488
rect 15151 3516 15163 3519
rect 17313 3519 17371 3525
rect 17313 3516 17325 3519
rect 15151 3488 17325 3516
rect 15151 3485 15163 3488
rect 15105 3479 15163 3485
rect 17313 3485 17325 3488
rect 17359 3485 17371 3519
rect 17313 3479 17371 3485
rect 17589 3519 17647 3525
rect 17589 3485 17601 3519
rect 17635 3516 17647 3519
rect 17678 3516 17684 3528
rect 17635 3488 17684 3516
rect 17635 3485 17647 3488
rect 17589 3479 17647 3485
rect 17678 3476 17684 3488
rect 17736 3476 17742 3528
rect 17954 3476 17960 3528
rect 18012 3516 18018 3528
rect 20346 3516 20352 3528
rect 18012 3488 20352 3516
rect 18012 3476 18018 3488
rect 16850 3448 16856 3460
rect 16811 3420 16856 3448
rect 16850 3408 16856 3420
rect 16908 3408 16914 3460
rect 19352 3448 19380 3488
rect 20346 3476 20352 3488
rect 20404 3516 20410 3528
rect 21836 3516 21864 3556
rect 22554 3544 22560 3556
rect 22612 3544 22618 3596
rect 25516 3593 25544 3624
rect 25774 3612 25780 3624
rect 25832 3612 25838 3664
rect 25866 3612 25872 3664
rect 25924 3652 25930 3664
rect 27154 3652 27160 3664
rect 25924 3624 25969 3652
rect 27115 3624 27160 3652
rect 25924 3612 25930 3624
rect 27154 3612 27160 3624
rect 27212 3612 27218 3664
rect 29638 3652 29644 3664
rect 28382 3624 29644 3652
rect 29638 3612 29644 3624
rect 29696 3612 29702 3664
rect 31772 3652 31800 3692
rect 36814 3680 36820 3692
rect 36872 3680 36878 3732
rect 36998 3680 37004 3732
rect 37056 3720 37062 3732
rect 37458 3720 37464 3732
rect 37056 3692 37320 3720
rect 37419 3692 37464 3720
rect 37056 3680 37062 3692
rect 31510 3624 31800 3652
rect 31846 3612 31852 3664
rect 31904 3652 31910 3664
rect 31904 3624 32260 3652
rect 31904 3612 31910 3624
rect 25501 3587 25559 3593
rect 20404 3488 21864 3516
rect 20404 3476 20410 3488
rect 19426 3448 19432 3460
rect 19352 3420 19432 3448
rect 19426 3408 19432 3420
rect 19484 3408 19490 3460
rect 23952 3448 23980 3570
rect 25501 3553 25513 3587
rect 25547 3553 25559 3587
rect 25501 3547 25559 3553
rect 24302 3516 24308 3528
rect 24263 3488 24308 3516
rect 24302 3476 24308 3488
rect 24360 3476 24366 3528
rect 25409 3519 25467 3525
rect 25409 3485 25421 3519
rect 25455 3516 25467 3519
rect 25884 3516 25912 3612
rect 26878 3584 26884 3596
rect 26839 3556 26884 3584
rect 26878 3544 26884 3556
rect 26936 3544 26942 3596
rect 28442 3544 28448 3596
rect 28500 3584 28506 3596
rect 29086 3584 29092 3596
rect 28500 3556 29092 3584
rect 28500 3544 28506 3556
rect 29086 3544 29092 3556
rect 29144 3544 29150 3596
rect 29273 3587 29331 3593
rect 29273 3553 29285 3587
rect 29319 3584 29331 3587
rect 29362 3584 29368 3596
rect 29319 3556 29368 3584
rect 29319 3553 29331 3556
rect 29273 3547 29331 3553
rect 29362 3544 29368 3556
rect 29420 3544 29426 3596
rect 31570 3516 31576 3528
rect 25455 3488 25912 3516
rect 26988 3488 31576 3516
rect 25455 3485 25467 3488
rect 25409 3479 25467 3485
rect 26988 3448 27016 3488
rect 31570 3476 31576 3488
rect 31628 3476 31634 3528
rect 31846 3476 31852 3528
rect 31904 3516 31910 3528
rect 32232 3525 32260 3624
rect 33134 3612 33140 3664
rect 33192 3612 33198 3664
rect 34146 3652 34152 3664
rect 34107 3624 34152 3652
rect 34146 3612 34152 3624
rect 34204 3612 34210 3664
rect 35986 3652 35992 3664
rect 35947 3624 35992 3652
rect 35986 3612 35992 3624
rect 36044 3612 36050 3664
rect 36446 3612 36452 3664
rect 36504 3612 36510 3664
rect 34425 3587 34483 3593
rect 34425 3553 34437 3587
rect 34471 3584 34483 3587
rect 34698 3584 34704 3596
rect 34471 3556 34704 3584
rect 34471 3553 34483 3556
rect 34425 3547 34483 3553
rect 31941 3519 31999 3525
rect 31941 3516 31953 3519
rect 31904 3488 31953 3516
rect 31904 3476 31910 3488
rect 31941 3485 31953 3488
rect 31987 3485 31999 3519
rect 31941 3479 31999 3485
rect 32217 3519 32275 3525
rect 32217 3485 32229 3519
rect 32263 3516 32275 3519
rect 33594 3516 33600 3528
rect 32263 3488 33600 3516
rect 32263 3485 32275 3488
rect 32217 3479 32275 3485
rect 33594 3476 33600 3488
rect 33652 3516 33658 3528
rect 34440 3516 34468 3547
rect 34698 3544 34704 3556
rect 34756 3584 34762 3596
rect 35713 3587 35771 3593
rect 35713 3584 35725 3587
rect 34756 3556 35725 3584
rect 34756 3544 34762 3556
rect 35713 3553 35725 3556
rect 35759 3553 35771 3587
rect 37292 3584 37320 3692
rect 37458 3680 37464 3692
rect 37516 3680 37522 3732
rect 37918 3720 37924 3732
rect 37879 3692 37924 3720
rect 37918 3680 37924 3692
rect 37976 3680 37982 3732
rect 38105 3587 38163 3593
rect 38105 3584 38117 3587
rect 37292 3556 38117 3584
rect 35713 3547 35771 3553
rect 38105 3553 38117 3556
rect 38151 3553 38163 3587
rect 38105 3547 38163 3553
rect 33652 3488 34468 3516
rect 33652 3476 33658 3488
rect 28718 3448 28724 3460
rect 23952 3420 27016 3448
rect 28460 3420 28724 3448
rect 17218 3340 17224 3392
rect 17276 3380 17282 3392
rect 22002 3380 22008 3392
rect 17276 3352 22008 3380
rect 17276 3340 17282 3352
rect 22002 3340 22008 3352
rect 22060 3340 22066 3392
rect 22097 3383 22155 3389
rect 22097 3349 22109 3383
rect 22143 3380 22155 3383
rect 23382 3380 23388 3392
rect 22143 3352 23388 3380
rect 22143 3349 22155 3352
rect 22097 3343 22155 3349
rect 23382 3340 23388 3352
rect 23440 3340 23446 3392
rect 24762 3340 24768 3392
rect 24820 3380 24826 3392
rect 28460 3380 28488 3420
rect 28718 3408 28724 3420
rect 28776 3408 28782 3460
rect 28810 3408 28816 3460
rect 28868 3448 28874 3460
rect 30469 3451 30527 3457
rect 30469 3448 30481 3451
rect 28868 3420 30481 3448
rect 28868 3408 28874 3420
rect 30469 3417 30481 3420
rect 30515 3417 30527 3451
rect 30469 3411 30527 3417
rect 24820 3352 28488 3380
rect 24820 3340 24826 3352
rect 28534 3340 28540 3392
rect 28592 3380 28598 3392
rect 29089 3383 29147 3389
rect 29089 3380 29101 3383
rect 28592 3352 29101 3380
rect 28592 3340 28598 3352
rect 29089 3349 29101 3352
rect 29135 3349 29147 3383
rect 29089 3343 29147 3349
rect 29178 3340 29184 3392
rect 29236 3380 29242 3392
rect 32306 3380 32312 3392
rect 29236 3352 32312 3380
rect 29236 3340 29242 3352
rect 32306 3340 32312 3352
rect 32364 3340 32370 3392
rect 32674 3380 32680 3392
rect 32635 3352 32680 3380
rect 32674 3340 32680 3352
rect 32732 3340 32738 3392
rect 32950 3340 32956 3392
rect 33008 3380 33014 3392
rect 34054 3380 34060 3392
rect 33008 3352 34060 3380
rect 33008 3340 33014 3352
rect 34054 3340 34060 3352
rect 34112 3380 34118 3392
rect 35434 3380 35440 3392
rect 34112 3352 35440 3380
rect 34112 3340 34118 3352
rect 35434 3340 35440 3352
rect 35492 3340 35498 3392
rect 1104 3290 38824 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 38824 3290
rect 1104 3216 38824 3238
rect 14093 3179 14151 3185
rect 14093 3145 14105 3179
rect 14139 3176 14151 3179
rect 17678 3176 17684 3188
rect 14139 3148 17540 3176
rect 17639 3148 17684 3176
rect 14139 3145 14151 3148
rect 14093 3139 14151 3145
rect 16393 3111 16451 3117
rect 16393 3077 16405 3111
rect 16439 3108 16451 3111
rect 16482 3108 16488 3120
rect 16439 3080 16488 3108
rect 16439 3077 16451 3080
rect 16393 3071 16451 3077
rect 16482 3068 16488 3080
rect 16540 3068 16546 3120
rect 17512 3108 17540 3148
rect 17678 3136 17684 3148
rect 17736 3136 17742 3188
rect 20152 3179 20210 3185
rect 20152 3145 20164 3179
rect 20198 3176 20210 3179
rect 21542 3176 21548 3188
rect 20198 3148 21548 3176
rect 20198 3145 20210 3148
rect 20152 3139 20210 3145
rect 21542 3136 21548 3148
rect 21600 3136 21606 3188
rect 21637 3179 21695 3185
rect 21637 3145 21649 3179
rect 21683 3176 21695 3179
rect 22830 3176 22836 3188
rect 21683 3148 22836 3176
rect 21683 3145 21695 3148
rect 21637 3139 21695 3145
rect 22830 3136 22836 3148
rect 22888 3136 22894 3188
rect 26881 3179 26939 3185
rect 26881 3145 26893 3179
rect 26927 3176 26939 3179
rect 27706 3176 27712 3188
rect 26927 3148 27712 3176
rect 26927 3145 26939 3148
rect 26881 3139 26939 3145
rect 27706 3136 27712 3148
rect 27764 3136 27770 3188
rect 29178 3176 29184 3188
rect 27908 3148 29184 3176
rect 23014 3108 23020 3120
rect 17512 3080 18184 3108
rect 18156 3040 18184 3080
rect 21192 3080 23020 3108
rect 21192 3040 21220 3080
rect 23014 3068 23020 3080
rect 23072 3068 23078 3120
rect 14200 3012 17908 3040
rect 18156 3012 21220 3040
rect 14200 2981 14228 3012
rect 14185 2975 14243 2981
rect 14185 2941 14197 2975
rect 14231 2941 14243 2975
rect 14642 2972 14648 2984
rect 14603 2944 14648 2972
rect 14185 2935 14243 2941
rect 14642 2932 14648 2944
rect 14700 2932 14706 2984
rect 14921 2907 14979 2913
rect 14921 2873 14933 2907
rect 14967 2904 14979 2907
rect 15194 2904 15200 2916
rect 14967 2876 15200 2904
rect 14967 2873 14979 2876
rect 14921 2867 14979 2873
rect 15194 2864 15200 2876
rect 15252 2864 15258 2916
rect 16482 2904 16488 2916
rect 16146 2876 16488 2904
rect 16482 2864 16488 2876
rect 16540 2864 16546 2916
rect 17880 2836 17908 3012
rect 21358 3000 21364 3052
rect 21416 3000 21422 3052
rect 21726 3000 21732 3052
rect 21784 3040 21790 3052
rect 22603 3043 22661 3049
rect 22603 3040 22615 3043
rect 21784 3012 22615 3040
rect 21784 3000 21790 3012
rect 22603 3009 22615 3012
rect 22649 3009 22661 3043
rect 24026 3040 24032 3052
rect 23987 3012 24032 3040
rect 22603 3003 22661 3009
rect 24026 3000 24032 3012
rect 24084 3000 24090 3052
rect 24397 3043 24455 3049
rect 24397 3009 24409 3043
rect 24443 3040 24455 3043
rect 25130 3040 25136 3052
rect 24443 3012 25136 3040
rect 24443 3009 24455 3012
rect 24397 3003 24455 3009
rect 25130 3000 25136 3012
rect 25188 3000 25194 3052
rect 25409 3043 25467 3049
rect 25409 3009 25421 3043
rect 25455 3040 25467 3043
rect 27522 3040 27528 3052
rect 25455 3012 27528 3040
rect 25455 3009 25467 3012
rect 25409 3003 25467 3009
rect 27522 3000 27528 3012
rect 27580 3000 27586 3052
rect 19426 2932 19432 2984
rect 19484 2972 19490 2984
rect 19886 2972 19892 2984
rect 19484 2944 19892 2972
rect 19484 2932 19490 2944
rect 19886 2932 19892 2944
rect 19944 2932 19950 2984
rect 21376 2972 21404 3000
rect 27908 2972 27936 3148
rect 29178 3136 29184 3148
rect 29236 3136 29242 3188
rect 30650 3136 30656 3188
rect 30708 3176 30714 3188
rect 31294 3176 31300 3188
rect 30708 3148 31300 3176
rect 30708 3136 30714 3148
rect 31294 3136 31300 3148
rect 31352 3136 31358 3188
rect 31570 3136 31576 3188
rect 31628 3176 31634 3188
rect 32674 3176 32680 3188
rect 31628 3148 32680 3176
rect 31628 3136 31634 3148
rect 32674 3136 32680 3148
rect 32732 3136 32738 3188
rect 33042 3176 33048 3188
rect 33003 3148 33048 3176
rect 33042 3136 33048 3148
rect 33100 3136 33106 3188
rect 34146 3136 34152 3188
rect 34204 3176 34210 3188
rect 36909 3179 36967 3185
rect 36909 3176 36921 3179
rect 34204 3148 36921 3176
rect 34204 3136 34210 3148
rect 36909 3145 36921 3148
rect 36955 3145 36967 3179
rect 36909 3139 36967 3145
rect 27982 3068 27988 3120
rect 28040 3108 28046 3120
rect 35253 3111 35311 3117
rect 28040 3080 28672 3108
rect 28040 3068 28046 3080
rect 28644 3049 28672 3080
rect 30392 3080 33548 3108
rect 28629 3043 28687 3049
rect 28629 3009 28641 3043
rect 28675 3009 28687 3043
rect 28629 3003 28687 3009
rect 28997 3043 29055 3049
rect 28997 3009 29009 3043
rect 29043 3040 29055 3043
rect 30392 3040 30420 3080
rect 29043 3012 30420 3040
rect 30929 3043 30987 3049
rect 29043 3009 29055 3012
rect 28997 3003 29055 3009
rect 30929 3009 30941 3043
rect 30975 3040 30987 3043
rect 31389 3043 31447 3049
rect 31389 3040 31401 3043
rect 30975 3012 31401 3040
rect 30975 3009 30987 3012
rect 30929 3003 30987 3009
rect 31389 3009 31401 3012
rect 31435 3009 31447 3043
rect 31389 3003 31447 3009
rect 21376 2944 23060 2972
rect 26542 2944 27936 2972
rect 27985 2975 28043 2981
rect 18690 2864 18696 2916
rect 18748 2864 18754 2916
rect 19058 2864 19064 2916
rect 19116 2904 19122 2916
rect 19153 2907 19211 2913
rect 19153 2904 19165 2907
rect 19116 2876 19165 2904
rect 19116 2864 19122 2876
rect 19153 2873 19165 2876
rect 19199 2873 19211 2907
rect 22002 2904 22008 2916
rect 21390 2876 22008 2904
rect 19153 2867 19211 2873
rect 22002 2864 22008 2876
rect 22060 2864 22066 2916
rect 23032 2890 23060 2944
rect 27985 2941 27997 2975
rect 28031 2972 28043 2975
rect 28534 2972 28540 2984
rect 28031 2944 28540 2972
rect 28031 2941 28043 2944
rect 27985 2935 28043 2941
rect 28534 2932 28540 2944
rect 28592 2932 28598 2984
rect 28902 2972 28908 2984
rect 28644 2944 28908 2972
rect 28644 2904 28672 2944
rect 28902 2932 28908 2944
rect 28960 2932 28966 2984
rect 31294 2972 31300 2984
rect 30024 2944 31156 2972
rect 31255 2944 31300 2972
rect 26712 2876 28672 2904
rect 30024 2890 30052 2944
rect 23934 2836 23940 2848
rect 17880 2808 23940 2836
rect 23934 2796 23940 2808
rect 23992 2836 23998 2848
rect 26712 2836 26740 2876
rect 30650 2864 30656 2916
rect 30708 2904 30714 2916
rect 31021 2907 31079 2913
rect 31021 2904 31033 2907
rect 30708 2876 31033 2904
rect 30708 2864 30714 2876
rect 31021 2873 31033 2876
rect 31067 2873 31079 2907
rect 31128 2904 31156 2944
rect 31294 2932 31300 2944
rect 31352 2932 31358 2984
rect 31404 2972 31432 3003
rect 31478 3000 31484 3052
rect 31536 3040 31542 3052
rect 33520 3040 33548 3080
rect 35253 3077 35265 3111
rect 35299 3077 35311 3111
rect 35253 3071 35311 3077
rect 35268 3040 35296 3071
rect 31536 3012 33088 3040
rect 33520 3012 35296 3040
rect 31536 3000 31542 3012
rect 32950 2972 32956 2984
rect 31404 2944 32956 2972
rect 32950 2932 32956 2944
rect 33008 2932 33014 2984
rect 32766 2904 32772 2916
rect 31128 2876 32772 2904
rect 31021 2867 31079 2873
rect 32766 2864 32772 2876
rect 32824 2864 32830 2916
rect 23992 2808 26740 2836
rect 28169 2839 28227 2845
rect 23992 2796 23998 2808
rect 28169 2805 28181 2839
rect 28215 2836 28227 2839
rect 30282 2836 30288 2848
rect 28215 2808 30288 2836
rect 28215 2805 28227 2808
rect 28169 2799 28227 2805
rect 30282 2796 30288 2808
rect 30340 2796 30346 2848
rect 30423 2839 30481 2845
rect 30423 2805 30435 2839
rect 30469 2836 30481 2839
rect 31478 2836 31484 2848
rect 30469 2808 31484 2836
rect 30469 2805 30481 2808
rect 30423 2799 30481 2805
rect 31478 2796 31484 2808
rect 31536 2796 31542 2848
rect 31573 2839 31631 2845
rect 31573 2805 31585 2839
rect 31619 2836 31631 2839
rect 32950 2836 32956 2848
rect 31619 2808 32956 2836
rect 31619 2805 31631 2808
rect 31573 2799 31631 2805
rect 32950 2796 32956 2808
rect 33008 2796 33014 2848
rect 33060 2836 33088 3012
rect 35342 3000 35348 3052
rect 35400 3040 35406 3052
rect 35400 3012 36400 3040
rect 35400 3000 35406 3012
rect 34790 2932 34796 2984
rect 34848 2972 34854 2984
rect 35434 2972 35440 2984
rect 34848 2944 34893 2972
rect 35395 2944 35440 2972
rect 34848 2932 34854 2944
rect 35434 2932 35440 2944
rect 35492 2932 35498 2984
rect 35526 2932 35532 2984
rect 35584 2972 35590 2984
rect 36372 2981 36400 3012
rect 36446 3000 36452 3052
rect 36504 3040 36510 3052
rect 36504 3012 36549 3040
rect 36504 3000 36510 3012
rect 35805 2975 35863 2981
rect 35805 2972 35817 2975
rect 35584 2944 35817 2972
rect 35584 2932 35590 2944
rect 35805 2941 35817 2944
rect 35851 2941 35863 2975
rect 35805 2935 35863 2941
rect 36357 2975 36415 2981
rect 36357 2941 36369 2975
rect 36403 2941 36415 2975
rect 36357 2935 36415 2941
rect 36633 2975 36691 2981
rect 36633 2941 36645 2975
rect 36679 2941 36691 2975
rect 36633 2935 36691 2941
rect 33134 2864 33140 2916
rect 33192 2904 33198 2916
rect 34514 2904 34520 2916
rect 33192 2876 33350 2904
rect 34475 2876 34520 2904
rect 33192 2864 33198 2876
rect 34514 2864 34520 2876
rect 34572 2864 34578 2916
rect 35452 2904 35480 2932
rect 35897 2907 35955 2913
rect 35897 2904 35909 2907
rect 35452 2876 35909 2904
rect 35897 2873 35909 2876
rect 35943 2904 35955 2907
rect 36648 2904 36676 2935
rect 36722 2932 36728 2984
rect 36780 2972 36786 2984
rect 36780 2944 36825 2972
rect 36780 2932 36786 2944
rect 35943 2876 36676 2904
rect 35943 2873 35955 2876
rect 35897 2867 35955 2873
rect 34606 2836 34612 2848
rect 33060 2808 34612 2836
rect 34606 2796 34612 2808
rect 34664 2796 34670 2848
rect 34698 2796 34704 2848
rect 34756 2836 34762 2848
rect 36446 2836 36452 2848
rect 34756 2808 36452 2836
rect 34756 2796 34762 2808
rect 36446 2796 36452 2808
rect 36504 2796 36510 2848
rect 1104 2746 38824 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 38824 2746
rect 1104 2672 38824 2694
rect 16022 2632 16028 2644
rect 15983 2604 16028 2632
rect 16022 2592 16028 2604
rect 16080 2592 16086 2644
rect 16482 2632 16488 2644
rect 16443 2604 16488 2632
rect 16482 2592 16488 2604
rect 16540 2592 16546 2644
rect 16574 2592 16580 2644
rect 16632 2632 16638 2644
rect 18230 2632 18236 2644
rect 16632 2604 18236 2632
rect 16632 2592 16638 2604
rect 18230 2592 18236 2604
rect 18288 2592 18294 2644
rect 19334 2632 19340 2644
rect 19295 2604 19340 2632
rect 19334 2592 19340 2604
rect 19392 2592 19398 2644
rect 21174 2632 21180 2644
rect 19720 2604 21180 2632
rect 15105 2567 15163 2573
rect 15105 2533 15117 2567
rect 15151 2564 15163 2567
rect 17402 2564 17408 2576
rect 15151 2536 17408 2564
rect 15151 2533 15163 2536
rect 15105 2527 15163 2533
rect 17402 2524 17408 2536
rect 17460 2524 17466 2576
rect 17862 2564 17868 2576
rect 17823 2536 17868 2564
rect 17862 2524 17868 2536
rect 17920 2524 17926 2576
rect 19720 2564 19748 2604
rect 21174 2592 21180 2604
rect 21232 2592 21238 2644
rect 22005 2635 22063 2641
rect 22005 2601 22017 2635
rect 22051 2632 22063 2635
rect 24118 2632 24124 2644
rect 22051 2604 24124 2632
rect 22051 2601 22063 2604
rect 22005 2595 22063 2601
rect 24118 2592 24124 2604
rect 24176 2592 24182 2644
rect 24673 2635 24731 2641
rect 24673 2601 24685 2635
rect 24719 2632 24731 2635
rect 24946 2632 24952 2644
rect 24719 2604 24952 2632
rect 24719 2601 24731 2604
rect 24673 2595 24731 2601
rect 24946 2592 24952 2604
rect 25004 2592 25010 2644
rect 26694 2592 26700 2644
rect 26752 2592 26758 2644
rect 27522 2592 27528 2644
rect 27580 2632 27586 2644
rect 30009 2635 30067 2641
rect 30009 2632 30021 2635
rect 27580 2604 30021 2632
rect 27580 2592 27586 2604
rect 30009 2601 30021 2604
rect 30055 2601 30067 2635
rect 30009 2595 30067 2601
rect 30929 2635 30987 2641
rect 30929 2601 30941 2635
rect 30975 2632 30987 2635
rect 31754 2632 31760 2644
rect 30975 2604 31760 2632
rect 30975 2601 30987 2604
rect 30929 2595 30987 2601
rect 31754 2592 31760 2604
rect 31812 2592 31818 2644
rect 34146 2632 34152 2644
rect 32416 2604 34152 2632
rect 19090 2536 19748 2564
rect 20990 2524 20996 2576
rect 21048 2524 21054 2576
rect 23201 2567 23259 2573
rect 23201 2533 23213 2567
rect 23247 2564 23259 2567
rect 23474 2564 23480 2576
rect 23247 2536 23480 2564
rect 23247 2533 23259 2536
rect 23201 2527 23259 2533
rect 23474 2524 23480 2536
rect 23532 2524 23538 2576
rect 26712 2564 26740 2592
rect 26634 2536 26740 2564
rect 27065 2567 27123 2573
rect 27065 2533 27077 2567
rect 27111 2564 27123 2567
rect 28810 2564 28816 2576
rect 27111 2536 28816 2564
rect 27111 2533 27123 2536
rect 27065 2527 27123 2533
rect 28810 2524 28816 2536
rect 28868 2524 28874 2576
rect 29914 2564 29920 2576
rect 29762 2536 29920 2564
rect 29914 2524 29920 2536
rect 29972 2524 29978 2576
rect 32416 2573 32444 2604
rect 34146 2592 34152 2604
rect 34204 2592 34210 2644
rect 35345 2635 35403 2641
rect 35345 2601 35357 2635
rect 35391 2632 35403 2635
rect 35526 2632 35532 2644
rect 35391 2604 35532 2632
rect 35391 2601 35403 2604
rect 35345 2595 35403 2601
rect 35526 2592 35532 2604
rect 35584 2592 35590 2644
rect 32401 2567 32459 2573
rect 32401 2533 32413 2567
rect 32447 2533 32459 2567
rect 32401 2527 32459 2533
rect 32950 2524 32956 2576
rect 33008 2564 33014 2576
rect 33873 2567 33931 2573
rect 33873 2564 33885 2567
rect 33008 2536 33885 2564
rect 33008 2524 33014 2536
rect 33873 2533 33885 2536
rect 33919 2533 33931 2567
rect 33873 2527 33931 2533
rect 34330 2524 34336 2576
rect 34388 2524 34394 2576
rect 36446 2564 36452 2576
rect 36407 2536 36452 2564
rect 36446 2524 36452 2536
rect 36504 2524 36510 2576
rect 13170 2496 13176 2508
rect 13131 2468 13176 2496
rect 13170 2456 13176 2468
rect 13228 2456 13234 2508
rect 13817 2499 13875 2505
rect 13817 2465 13829 2499
rect 13863 2496 13875 2499
rect 15841 2499 15899 2505
rect 15841 2496 15853 2499
rect 13863 2468 15853 2496
rect 13863 2465 13875 2468
rect 13817 2459 13875 2465
rect 15841 2465 15853 2468
rect 15887 2496 15899 2499
rect 16669 2499 16727 2505
rect 15887 2468 16574 2496
rect 15887 2465 15899 2468
rect 15841 2459 15899 2465
rect 16546 2440 16574 2468
rect 16669 2465 16681 2499
rect 16715 2465 16727 2499
rect 16669 2459 16727 2465
rect 16546 2400 16580 2440
rect 16574 2388 16580 2400
rect 16632 2388 16638 2440
rect 14918 2360 14924 2372
rect 14879 2332 14924 2360
rect 14918 2320 14924 2332
rect 14976 2320 14982 2372
rect 13354 2292 13360 2304
rect 13315 2264 13360 2292
rect 13354 2252 13360 2264
rect 13412 2252 13418 2304
rect 13998 2292 14004 2304
rect 13959 2264 14004 2292
rect 13998 2252 14004 2264
rect 14056 2252 14062 2304
rect 16684 2292 16712 2459
rect 19886 2456 19892 2508
rect 19944 2496 19950 2508
rect 20257 2499 20315 2505
rect 20257 2496 20269 2499
rect 19944 2468 20269 2496
rect 19944 2456 19950 2468
rect 20257 2465 20269 2468
rect 20303 2465 20315 2499
rect 20257 2459 20315 2465
rect 22554 2456 22560 2508
rect 22612 2496 22618 2508
rect 22925 2499 22983 2505
rect 22925 2496 22937 2499
rect 22612 2468 22937 2496
rect 22612 2456 22618 2468
rect 22925 2465 22937 2468
rect 22971 2465 22983 2499
rect 22925 2459 22983 2465
rect 24302 2456 24308 2508
rect 24360 2456 24366 2508
rect 27341 2499 27399 2505
rect 27341 2465 27353 2499
rect 27387 2496 27399 2499
rect 27798 2496 27804 2508
rect 27387 2468 27804 2496
rect 27387 2465 27399 2468
rect 27341 2459 27399 2465
rect 27798 2456 27804 2468
rect 27856 2496 27862 2508
rect 28261 2499 28319 2505
rect 28261 2496 28273 2499
rect 27856 2468 28273 2496
rect 27856 2456 27862 2468
rect 28261 2465 28273 2468
rect 28307 2465 28319 2499
rect 32677 2499 32735 2505
rect 28261 2459 28319 2465
rect 17494 2388 17500 2440
rect 17552 2428 17558 2440
rect 17589 2431 17647 2437
rect 17589 2428 17601 2431
rect 17552 2400 17601 2428
rect 17552 2388 17558 2400
rect 17589 2397 17601 2400
rect 17635 2397 17647 2431
rect 20530 2428 20536 2440
rect 20491 2400 20536 2428
rect 17589 2391 17647 2397
rect 20530 2388 20536 2400
rect 20588 2388 20594 2440
rect 24854 2388 24860 2440
rect 24912 2428 24918 2440
rect 25593 2431 25651 2437
rect 25593 2428 25605 2431
rect 24912 2400 25605 2428
rect 24912 2388 24918 2400
rect 25593 2397 25605 2400
rect 25639 2397 25651 2431
rect 25593 2391 25651 2397
rect 25682 2388 25688 2440
rect 25740 2428 25746 2440
rect 28537 2431 28595 2437
rect 28537 2428 28549 2431
rect 25740 2400 27292 2428
rect 25740 2388 25746 2400
rect 27264 2360 27292 2400
rect 28368 2400 28549 2428
rect 28368 2360 28396 2400
rect 28537 2397 28549 2400
rect 28583 2397 28595 2431
rect 31312 2428 31340 2482
rect 32677 2465 32689 2499
rect 32723 2496 32735 2499
rect 33594 2496 33600 2508
rect 32723 2468 33600 2496
rect 32723 2465 32735 2468
rect 32677 2459 32735 2465
rect 33594 2456 33600 2468
rect 33652 2456 33658 2508
rect 36906 2456 36912 2508
rect 36964 2496 36970 2508
rect 37185 2499 37243 2505
rect 37185 2496 37197 2499
rect 36964 2468 37197 2496
rect 36964 2456 36970 2468
rect 37185 2465 37197 2468
rect 37231 2465 37243 2499
rect 37826 2496 37832 2508
rect 37787 2468 37832 2496
rect 37185 2459 37243 2465
rect 37826 2456 37832 2468
rect 37884 2456 37890 2508
rect 31312 2400 32628 2428
rect 28537 2391 28595 2397
rect 27264 2332 28396 2360
rect 32600 2360 32628 2400
rect 32858 2388 32864 2440
rect 32916 2428 32922 2440
rect 32916 2400 37688 2428
rect 32916 2388 32922 2400
rect 33502 2360 33508 2372
rect 32600 2332 33508 2360
rect 33502 2320 33508 2332
rect 33560 2320 33566 2372
rect 35250 2320 35256 2372
rect 35308 2360 35314 2372
rect 37660 2369 37688 2400
rect 36265 2363 36323 2369
rect 36265 2360 36277 2363
rect 35308 2332 36277 2360
rect 35308 2320 35314 2332
rect 36265 2329 36277 2332
rect 36311 2329 36323 2363
rect 36265 2323 36323 2329
rect 37645 2363 37703 2369
rect 37645 2329 37657 2363
rect 37691 2329 37703 2363
rect 37645 2323 37703 2329
rect 25222 2292 25228 2304
rect 16684 2264 25228 2292
rect 25222 2252 25228 2264
rect 25280 2252 25286 2304
rect 36998 2292 37004 2304
rect 36959 2264 37004 2292
rect 36998 2252 37004 2264
rect 37056 2252 37062 2304
rect 1104 2202 38824 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 38824 2202
rect 1104 2128 38824 2150
rect 13354 2048 13360 2100
rect 13412 2088 13418 2100
rect 20530 2088 20536 2100
rect 13412 2060 20536 2088
rect 13412 2048 13418 2060
rect 20530 2048 20536 2060
rect 20588 2048 20594 2100
rect 22002 2048 22008 2100
rect 22060 2088 22066 2100
rect 36998 2088 37004 2100
rect 22060 2060 37004 2088
rect 22060 2048 22066 2060
rect 36998 2048 37004 2060
rect 37056 2048 37062 2100
rect 13998 1980 14004 2032
rect 14056 2020 14062 2032
rect 20990 2020 20996 2032
rect 14056 1992 20996 2020
rect 14056 1980 14062 1992
rect 20990 1980 20996 1992
rect 21048 1980 21054 2032
rect 24302 1980 24308 2032
rect 24360 2020 24366 2032
rect 24360 1992 26234 2020
rect 24360 1980 24366 1992
rect 13170 1912 13176 1964
rect 13228 1952 13234 1964
rect 24946 1952 24952 1964
rect 13228 1924 24952 1952
rect 13228 1912 13234 1924
rect 24946 1912 24952 1924
rect 25004 1912 25010 1964
rect 26206 1952 26234 1992
rect 29086 1980 29092 2032
rect 29144 2020 29150 2032
rect 34330 2020 34336 2032
rect 29144 1992 34336 2020
rect 29144 1980 29150 1992
rect 34330 1980 34336 1992
rect 34388 1980 34394 2032
rect 31110 1952 31116 1964
rect 26206 1924 31116 1952
rect 31110 1912 31116 1924
rect 31168 1912 31174 1964
<< via1 >>
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 38108 19907 38160 19916
rect 38108 19873 38117 19907
rect 38117 19873 38151 19907
rect 38151 19873 38160 19907
rect 38108 19864 38160 19873
rect 35256 19660 35308 19712
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 35256 13472 35308 13524
rect 33048 13404 33100 13456
rect 33416 13311 33468 13320
rect 33416 13277 33425 13311
rect 33425 13277 33459 13311
rect 33459 13277 33468 13311
rect 33416 13268 33468 13277
rect 32220 13132 32272 13184
rect 32956 13132 33008 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 33416 12928 33468 12980
rect 31852 12792 31904 12844
rect 30656 12767 30708 12776
rect 30656 12733 30665 12767
rect 30665 12733 30699 12767
rect 30699 12733 30708 12767
rect 30656 12724 30708 12733
rect 32956 12724 33008 12776
rect 35256 12656 35308 12708
rect 32680 12588 32732 12640
rect 33048 12588 33100 12640
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 33048 12316 33100 12368
rect 30656 12248 30708 12300
rect 32220 12291 32272 12300
rect 32220 12257 32229 12291
rect 32229 12257 32263 12291
rect 32263 12257 32272 12291
rect 32220 12248 32272 12257
rect 31852 12223 31904 12232
rect 31852 12189 31861 12223
rect 31861 12189 31895 12223
rect 31895 12189 31904 12223
rect 31852 12180 31904 12189
rect 33048 12044 33100 12096
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 32680 11228 32732 11280
rect 27712 11160 27764 11212
rect 33048 11203 33100 11212
rect 33048 11169 33057 11203
rect 33057 11169 33091 11203
rect 33091 11169 33100 11203
rect 33048 11160 33100 11169
rect 31852 11092 31904 11144
rect 23664 11024 23716 11076
rect 31392 11024 31444 11076
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 24124 10684 24176 10736
rect 27252 10616 27304 10668
rect 27896 10548 27948 10600
rect 30840 10548 30892 10600
rect 31024 10480 31076 10532
rect 27804 10455 27856 10464
rect 27804 10421 27813 10455
rect 27813 10421 27847 10455
rect 27847 10421 27856 10455
rect 27804 10412 27856 10421
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 31852 10208 31904 10260
rect 22836 10072 22888 10124
rect 25872 10072 25924 10124
rect 28908 10140 28960 10192
rect 27712 10115 27764 10124
rect 27712 10081 27721 10115
rect 27721 10081 27755 10115
rect 27755 10081 27764 10115
rect 27712 10072 27764 10081
rect 30840 10115 30892 10124
rect 28080 10004 28132 10056
rect 29920 10004 29972 10056
rect 30840 10081 30849 10115
rect 30849 10081 30883 10115
rect 30883 10081 30892 10115
rect 30840 10072 30892 10081
rect 31208 10004 31260 10056
rect 24952 9936 25004 9988
rect 26700 9936 26752 9988
rect 24308 9911 24360 9920
rect 24308 9877 24317 9911
rect 24317 9877 24351 9911
rect 24351 9877 24360 9911
rect 24308 9868 24360 9877
rect 25780 9911 25832 9920
rect 25780 9877 25789 9911
rect 25789 9877 25823 9911
rect 25823 9877 25832 9911
rect 25780 9868 25832 9877
rect 26332 9868 26384 9920
rect 29092 9868 29144 9920
rect 30656 9868 30708 9920
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 16120 9664 16172 9716
rect 25780 9664 25832 9716
rect 23112 9596 23164 9648
rect 28724 9596 28776 9648
rect 27528 9528 27580 9580
rect 22928 9460 22980 9512
rect 24676 9503 24728 9512
rect 24676 9469 24685 9503
rect 24685 9469 24719 9503
rect 24719 9469 24728 9503
rect 24676 9460 24728 9469
rect 25872 9460 25924 9512
rect 27620 9460 27672 9512
rect 28908 9460 28960 9512
rect 29092 9460 29144 9512
rect 4988 9392 5040 9444
rect 27436 9392 27488 9444
rect 29920 9503 29972 9512
rect 29920 9469 29937 9503
rect 29937 9469 29971 9503
rect 29971 9469 29972 9503
rect 32036 9528 32088 9580
rect 29920 9460 29972 9469
rect 31668 9460 31720 9512
rect 21272 9324 21324 9376
rect 25412 9324 25464 9376
rect 27252 9324 27304 9376
rect 28540 9324 28592 9376
rect 30472 9392 30524 9444
rect 29184 9324 29236 9376
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 22376 9120 22428 9172
rect 22836 9163 22888 9172
rect 22836 9129 22845 9163
rect 22845 9129 22879 9163
rect 22879 9129 22888 9163
rect 22836 9120 22888 9129
rect 20720 8984 20772 9036
rect 25412 9052 25464 9104
rect 26240 9052 26292 9104
rect 30288 9052 30340 9104
rect 23664 9027 23716 9036
rect 23664 8993 23673 9027
rect 23673 8993 23707 9027
rect 23707 8993 23716 9027
rect 23664 8984 23716 8993
rect 23848 8916 23900 8968
rect 27620 8984 27672 9036
rect 28080 9027 28132 9036
rect 28080 8993 28089 9027
rect 28089 8993 28123 9027
rect 28123 8993 28132 9027
rect 28080 8984 28132 8993
rect 28908 9027 28960 9036
rect 28908 8993 28917 9027
rect 28917 8993 28951 9027
rect 28951 8993 28960 9027
rect 28908 8984 28960 8993
rect 29092 8984 29144 9036
rect 30196 8984 30248 9036
rect 30656 9027 30708 9036
rect 30656 8993 30665 9027
rect 30665 8993 30699 9027
rect 30699 8993 30708 9027
rect 30656 8984 30708 8993
rect 37832 8984 37884 9036
rect 27804 8916 27856 8968
rect 27896 8916 27948 8968
rect 30104 8916 30156 8968
rect 27252 8848 27304 8900
rect 30472 8891 30524 8900
rect 23664 8780 23716 8832
rect 24768 8780 24820 8832
rect 25044 8780 25096 8832
rect 28080 8780 28132 8832
rect 28172 8780 28224 8832
rect 28908 8780 28960 8832
rect 30472 8857 30481 8891
rect 30481 8857 30515 8891
rect 30515 8857 30524 8891
rect 30472 8848 30524 8857
rect 30380 8780 30432 8832
rect 31484 8916 31536 8968
rect 30840 8848 30892 8900
rect 35440 8780 35492 8832
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 27712 8576 27764 8628
rect 20444 8508 20496 8560
rect 24308 8508 24360 8560
rect 28816 8440 28868 8492
rect 29184 8440 29236 8492
rect 30104 8576 30156 8628
rect 31208 8576 31260 8628
rect 29552 8508 29604 8560
rect 22928 8372 22980 8424
rect 22008 8304 22060 8356
rect 23848 8372 23900 8424
rect 23020 8279 23072 8288
rect 23020 8245 23029 8279
rect 23029 8245 23063 8279
rect 23063 8245 23072 8279
rect 23020 8236 23072 8245
rect 23480 8279 23532 8288
rect 23480 8245 23489 8279
rect 23489 8245 23523 8279
rect 23523 8245 23532 8279
rect 23480 8236 23532 8245
rect 29552 8415 29604 8424
rect 29552 8381 29561 8415
rect 29561 8381 29595 8415
rect 29595 8381 29604 8415
rect 32680 8440 32732 8492
rect 29552 8372 29604 8381
rect 31392 8415 31444 8424
rect 31392 8381 31401 8415
rect 31401 8381 31435 8415
rect 31435 8381 31444 8415
rect 31392 8372 31444 8381
rect 31668 8372 31720 8424
rect 24400 8304 24452 8356
rect 27896 8304 27948 8356
rect 24676 8236 24728 8288
rect 25228 8236 25280 8288
rect 27804 8279 27856 8288
rect 27804 8245 27813 8279
rect 27813 8245 27847 8279
rect 27847 8245 27856 8279
rect 27804 8236 27856 8245
rect 35716 8304 35768 8356
rect 31484 8236 31536 8288
rect 33140 8236 33192 8288
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 18972 8032 19024 8084
rect 19432 7964 19484 8016
rect 21548 7896 21600 7948
rect 22376 7828 22428 7880
rect 22468 7760 22520 7812
rect 18236 7692 18288 7744
rect 21548 7692 21600 7744
rect 21916 7735 21968 7744
rect 21916 7701 21925 7735
rect 21925 7701 21959 7735
rect 21959 7701 21968 7735
rect 21916 7692 21968 7701
rect 23020 7964 23072 8016
rect 36544 8032 36596 8084
rect 27804 7964 27856 8016
rect 28632 7964 28684 8016
rect 24308 7939 24360 7948
rect 24308 7905 24317 7939
rect 24317 7905 24351 7939
rect 24351 7905 24360 7939
rect 24308 7896 24360 7905
rect 25504 7871 25556 7880
rect 23572 7692 23624 7744
rect 25504 7837 25513 7871
rect 25513 7837 25547 7871
rect 25547 7837 25556 7871
rect 25504 7828 25556 7837
rect 27712 7828 27764 7880
rect 28080 7828 28132 7880
rect 32496 7964 32548 8016
rect 30656 7939 30708 7948
rect 30656 7905 30665 7939
rect 30665 7905 30699 7939
rect 30699 7905 30708 7939
rect 30656 7896 30708 7905
rect 30196 7828 30248 7880
rect 32036 7896 32088 7948
rect 33140 7896 33192 7948
rect 34612 7896 34664 7948
rect 31576 7828 31628 7880
rect 30840 7760 30892 7812
rect 30932 7760 30984 7812
rect 26976 7735 27028 7744
rect 26976 7701 26985 7735
rect 26985 7701 27019 7735
rect 27019 7701 27028 7735
rect 26976 7692 27028 7701
rect 27896 7692 27948 7744
rect 31116 7735 31168 7744
rect 31116 7701 31125 7735
rect 31125 7701 31159 7735
rect 31159 7701 31168 7735
rect 31116 7692 31168 7701
rect 31852 7692 31904 7744
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 21456 7420 21508 7472
rect 17868 7352 17920 7404
rect 25412 7488 25464 7540
rect 26240 7488 26292 7540
rect 30748 7488 30800 7540
rect 29920 7420 29972 7472
rect 30932 7420 30984 7472
rect 20628 7284 20680 7336
rect 21364 7284 21416 7336
rect 22100 7284 22152 7336
rect 22928 7284 22980 7336
rect 23020 7284 23072 7336
rect 24308 7352 24360 7404
rect 24584 7395 24636 7404
rect 24584 7361 24593 7395
rect 24593 7361 24627 7395
rect 24627 7361 24636 7395
rect 24584 7352 24636 7361
rect 28632 7352 28684 7404
rect 23940 7284 23992 7336
rect 29552 7327 29604 7336
rect 29552 7293 29561 7327
rect 29561 7293 29595 7327
rect 29595 7293 29604 7327
rect 30196 7352 30248 7404
rect 29552 7284 29604 7293
rect 30840 7327 30892 7336
rect 30840 7293 30849 7327
rect 30849 7293 30883 7327
rect 30883 7293 30892 7327
rect 30840 7284 30892 7293
rect 30932 7284 30984 7336
rect 31392 7284 31444 7336
rect 36912 7352 36964 7404
rect 33140 7284 33192 7336
rect 16028 7216 16080 7268
rect 24860 7259 24912 7268
rect 20076 7191 20128 7200
rect 20076 7157 20085 7191
rect 20085 7157 20119 7191
rect 20119 7157 20128 7191
rect 20076 7148 20128 7157
rect 21824 7148 21876 7200
rect 24860 7225 24869 7259
rect 24869 7225 24903 7259
rect 24903 7225 24912 7259
rect 24860 7216 24912 7225
rect 28540 7216 28592 7268
rect 25780 7148 25832 7200
rect 26424 7148 26476 7200
rect 27896 7148 27948 7200
rect 32956 7216 33008 7268
rect 33692 7284 33744 7336
rect 34152 7216 34204 7268
rect 30196 7191 30248 7200
rect 30196 7157 30205 7191
rect 30205 7157 30239 7191
rect 30239 7157 30248 7191
rect 30196 7148 30248 7157
rect 30656 7148 30708 7200
rect 30932 7148 30984 7200
rect 31300 7191 31352 7200
rect 31300 7157 31309 7191
rect 31309 7157 31343 7191
rect 31343 7157 31352 7191
rect 31300 7148 31352 7157
rect 31944 7148 31996 7200
rect 34060 7148 34112 7200
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 23112 6876 23164 6928
rect 28172 6944 28224 6996
rect 30012 6944 30064 6996
rect 31576 6944 31628 6996
rect 32036 6944 32088 6996
rect 34704 6944 34756 6996
rect 19892 6740 19944 6792
rect 16488 6672 16540 6724
rect 22560 6783 22612 6792
rect 22560 6749 22569 6783
rect 22569 6749 22603 6783
rect 22603 6749 22612 6783
rect 22560 6740 22612 6749
rect 26424 6876 26476 6928
rect 28908 6876 28960 6928
rect 30196 6876 30248 6928
rect 31668 6876 31720 6928
rect 24216 6808 24268 6860
rect 24400 6740 24452 6792
rect 28540 6808 28592 6860
rect 27344 6740 27396 6792
rect 27804 6783 27856 6792
rect 27804 6749 27813 6783
rect 27813 6749 27847 6783
rect 27847 6749 27856 6783
rect 27804 6740 27856 6749
rect 25228 6672 25280 6724
rect 22192 6604 22244 6656
rect 22928 6604 22980 6656
rect 27344 6604 27396 6656
rect 27620 6604 27672 6656
rect 27712 6604 27764 6656
rect 29552 6808 29604 6860
rect 32312 6808 32364 6860
rect 32680 6851 32732 6860
rect 31484 6740 31536 6792
rect 31576 6740 31628 6792
rect 31852 6740 31904 6792
rect 32404 6740 32456 6792
rect 32680 6817 32689 6851
rect 32689 6817 32723 6851
rect 32723 6817 32732 6851
rect 32680 6808 32732 6817
rect 33048 6808 33100 6860
rect 33416 6808 33468 6860
rect 34152 6851 34204 6860
rect 34152 6817 34161 6851
rect 34161 6817 34195 6851
rect 34195 6817 34204 6851
rect 34152 6808 34204 6817
rect 34612 6851 34664 6860
rect 34612 6817 34621 6851
rect 34621 6817 34655 6851
rect 34655 6817 34664 6851
rect 34612 6808 34664 6817
rect 35808 6808 35860 6860
rect 35900 6740 35952 6792
rect 33140 6672 33192 6724
rect 29276 6604 29328 6656
rect 30656 6604 30708 6656
rect 31760 6604 31812 6656
rect 32772 6604 32824 6656
rect 34612 6604 34664 6656
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 20260 6400 20312 6452
rect 22376 6400 22428 6452
rect 18880 6196 18932 6248
rect 22100 6264 22152 6316
rect 19892 6239 19944 6248
rect 19892 6205 19901 6239
rect 19901 6205 19935 6239
rect 19935 6205 19944 6239
rect 19892 6196 19944 6205
rect 22560 6264 22612 6316
rect 24492 6332 24544 6384
rect 25504 6400 25556 6452
rect 24952 6332 25004 6384
rect 27620 6332 27672 6384
rect 30472 6332 30524 6384
rect 31852 6400 31904 6452
rect 32220 6400 32272 6452
rect 32312 6400 32364 6452
rect 28080 6264 28132 6316
rect 29460 6264 29512 6316
rect 30748 6264 30800 6316
rect 31852 6264 31904 6316
rect 32036 6332 32088 6384
rect 34336 6264 34388 6316
rect 24584 6196 24636 6248
rect 27712 6196 27764 6248
rect 32128 6196 32180 6248
rect 19064 6128 19116 6180
rect 22100 6128 22152 6180
rect 24952 6128 25004 6180
rect 27436 6128 27488 6180
rect 28080 6171 28132 6180
rect 28080 6137 28089 6171
rect 28089 6137 28123 6171
rect 28123 6137 28132 6171
rect 28080 6128 28132 6137
rect 30196 6128 30248 6180
rect 31024 6128 31076 6180
rect 31484 6171 31536 6180
rect 31484 6137 31493 6171
rect 31493 6137 31527 6171
rect 31527 6137 31536 6171
rect 31484 6128 31536 6137
rect 32956 6196 33008 6248
rect 33876 6239 33928 6248
rect 33876 6205 33885 6239
rect 33885 6205 33919 6239
rect 33919 6205 33928 6239
rect 33876 6196 33928 6205
rect 34704 6264 34756 6316
rect 35532 6264 35584 6316
rect 35348 6196 35400 6248
rect 36084 6128 36136 6180
rect 18696 6060 18748 6112
rect 28816 6060 28868 6112
rect 30104 6060 30156 6112
rect 36728 6060 36780 6112
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 21364 5856 21416 5908
rect 15568 5720 15620 5772
rect 20076 5788 20128 5840
rect 24124 5788 24176 5840
rect 24860 5856 24912 5908
rect 30104 5856 30156 5908
rect 30288 5856 30340 5908
rect 31576 5856 31628 5908
rect 33048 5856 33100 5908
rect 35716 5899 35768 5908
rect 35716 5865 35725 5899
rect 35725 5865 35759 5899
rect 35759 5865 35768 5899
rect 35716 5856 35768 5865
rect 31852 5788 31904 5840
rect 18236 5763 18288 5772
rect 18236 5729 18245 5763
rect 18245 5729 18279 5763
rect 18279 5729 18288 5763
rect 18236 5720 18288 5729
rect 20260 5720 20312 5772
rect 22560 5763 22612 5772
rect 22560 5729 22569 5763
rect 22569 5729 22603 5763
rect 22603 5729 22612 5763
rect 22560 5720 22612 5729
rect 19892 5652 19944 5704
rect 20628 5695 20680 5704
rect 20628 5661 20637 5695
rect 20637 5661 20671 5695
rect 20671 5661 20680 5695
rect 20628 5652 20680 5661
rect 21640 5584 21692 5636
rect 23388 5652 23440 5704
rect 27160 5720 27212 5772
rect 29000 5720 29052 5772
rect 30380 5720 30432 5772
rect 25412 5695 25464 5704
rect 25412 5661 25421 5695
rect 25421 5661 25455 5695
rect 25455 5661 25464 5695
rect 25872 5695 25924 5704
rect 25412 5652 25464 5661
rect 25872 5661 25881 5695
rect 25881 5661 25915 5695
rect 25915 5661 25924 5695
rect 25872 5652 25924 5661
rect 24308 5584 24360 5636
rect 28080 5652 28132 5704
rect 28448 5695 28500 5704
rect 28448 5661 28457 5695
rect 28457 5661 28491 5695
rect 28491 5661 28500 5695
rect 28448 5652 28500 5661
rect 27436 5584 27488 5636
rect 28816 5652 28868 5704
rect 32220 5695 32272 5704
rect 32220 5661 32229 5695
rect 32229 5661 32263 5695
rect 32263 5661 32272 5695
rect 32220 5652 32272 5661
rect 32772 5788 32824 5840
rect 33876 5788 33928 5840
rect 32864 5763 32916 5772
rect 32864 5729 32873 5763
rect 32873 5729 32907 5763
rect 32907 5729 32916 5763
rect 32864 5720 32916 5729
rect 32956 5720 33008 5772
rect 35900 5763 35952 5772
rect 35900 5729 35909 5763
rect 35909 5729 35943 5763
rect 35943 5729 35952 5763
rect 35900 5720 35952 5729
rect 36820 5652 36872 5704
rect 17500 5516 17552 5568
rect 18880 5559 18932 5568
rect 18880 5525 18889 5559
rect 18889 5525 18923 5559
rect 18923 5525 18932 5559
rect 18880 5516 18932 5525
rect 21180 5516 21232 5568
rect 24032 5516 24084 5568
rect 27804 5516 27856 5568
rect 27988 5516 28040 5568
rect 30012 5584 30064 5636
rect 30196 5584 30248 5636
rect 29368 5559 29420 5568
rect 29368 5525 29377 5559
rect 29377 5525 29411 5559
rect 29411 5525 29420 5559
rect 29368 5516 29420 5525
rect 29828 5516 29880 5568
rect 32772 5516 32824 5568
rect 33324 5559 33376 5568
rect 33324 5525 33333 5559
rect 33333 5525 33367 5559
rect 33367 5525 33376 5559
rect 33324 5516 33376 5525
rect 33416 5516 33468 5568
rect 36452 5516 36504 5568
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 17316 5312 17368 5364
rect 19340 5312 19392 5364
rect 21732 5312 21784 5364
rect 23112 5312 23164 5364
rect 35716 5312 35768 5364
rect 17500 5176 17552 5228
rect 19892 5219 19944 5228
rect 19892 5185 19901 5219
rect 19901 5185 19935 5219
rect 19935 5185 19944 5219
rect 19892 5176 19944 5185
rect 21180 5176 21232 5228
rect 22836 5176 22888 5228
rect 25136 5244 25188 5296
rect 22468 5108 22520 5160
rect 27436 5176 27488 5228
rect 28816 5176 28868 5228
rect 29644 5244 29696 5296
rect 29552 5219 29604 5228
rect 29552 5185 29561 5219
rect 29561 5185 29595 5219
rect 29595 5185 29604 5219
rect 29552 5176 29604 5185
rect 29736 5176 29788 5228
rect 33048 5244 33100 5296
rect 35992 5244 36044 5296
rect 25136 5151 25188 5160
rect 25136 5117 25145 5151
rect 25145 5117 25179 5151
rect 25179 5117 25188 5151
rect 25136 5108 25188 5117
rect 20444 5040 20496 5092
rect 15200 4972 15252 5024
rect 19984 4972 20036 5024
rect 22836 5040 22888 5092
rect 23664 5040 23716 5092
rect 24124 5040 24176 5092
rect 25412 5083 25464 5092
rect 25412 5049 25421 5083
rect 25421 5049 25455 5083
rect 25455 5049 25464 5083
rect 25412 5040 25464 5049
rect 27528 5040 27580 5092
rect 21548 4972 21600 5024
rect 25504 4972 25556 5024
rect 27712 4972 27764 5024
rect 29000 5040 29052 5092
rect 30380 5040 30432 5092
rect 30564 5040 30616 5092
rect 31300 5040 31352 5092
rect 32220 5108 32272 5160
rect 33048 5151 33100 5160
rect 33048 5117 33057 5151
rect 33057 5117 33091 5151
rect 33091 5117 33100 5151
rect 33048 5108 33100 5117
rect 35440 5151 35492 5160
rect 35440 5117 35449 5151
rect 35449 5117 35483 5151
rect 35483 5117 35492 5151
rect 35440 5108 35492 5117
rect 35532 5108 35584 5160
rect 32496 5040 32548 5092
rect 33784 5040 33836 5092
rect 35900 5040 35952 5092
rect 32220 4972 32272 5024
rect 34244 4972 34296 5024
rect 34336 4972 34388 5024
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 18880 4768 18932 4820
rect 19340 4768 19392 4820
rect 21456 4768 21508 4820
rect 17500 4700 17552 4752
rect 35808 4768 35860 4820
rect 17592 4607 17644 4616
rect 17592 4573 17601 4607
rect 17601 4573 17635 4607
rect 17635 4573 17644 4607
rect 17592 4564 17644 4573
rect 18052 4428 18104 4480
rect 19156 4428 19208 4480
rect 20352 4607 20404 4616
rect 20352 4573 20361 4607
rect 20361 4573 20395 4607
rect 20395 4573 20404 4607
rect 20352 4564 20404 4573
rect 23112 4700 23164 4752
rect 25504 4743 25556 4752
rect 25504 4709 25513 4743
rect 25513 4709 25547 4743
rect 25547 4709 25556 4743
rect 25504 4700 25556 4709
rect 27436 4700 27488 4752
rect 27712 4743 27764 4752
rect 27712 4709 27721 4743
rect 27721 4709 27755 4743
rect 27755 4709 27764 4743
rect 27712 4700 27764 4709
rect 28356 4700 28408 4752
rect 30012 4700 30064 4752
rect 30748 4743 30800 4752
rect 22100 4607 22152 4616
rect 22100 4573 22109 4607
rect 22109 4573 22143 4607
rect 22143 4573 22152 4607
rect 22560 4607 22612 4616
rect 22100 4564 22152 4573
rect 22560 4573 22569 4607
rect 22569 4573 22603 4607
rect 22603 4573 22612 4607
rect 22560 4564 22612 4573
rect 22836 4607 22888 4616
rect 22836 4573 22845 4607
rect 22845 4573 22879 4607
rect 22879 4573 22888 4607
rect 22836 4564 22888 4573
rect 23204 4564 23256 4616
rect 23480 4564 23532 4616
rect 25136 4632 25188 4684
rect 27436 4607 27488 4616
rect 27436 4573 27445 4607
rect 27445 4573 27479 4607
rect 27479 4573 27488 4607
rect 27436 4564 27488 4573
rect 30380 4632 30432 4684
rect 30748 4709 30757 4743
rect 30757 4709 30791 4743
rect 30791 4709 30800 4743
rect 30748 4700 30800 4709
rect 32864 4700 32916 4752
rect 35256 4700 35308 4752
rect 34520 4632 34572 4684
rect 35348 4632 35400 4684
rect 35440 4632 35492 4684
rect 36360 4632 36412 4684
rect 36820 4632 36872 4684
rect 37832 4675 37884 4684
rect 29184 4607 29236 4616
rect 29184 4573 29193 4607
rect 29193 4573 29227 4607
rect 29227 4573 29236 4607
rect 29184 4564 29236 4573
rect 31484 4564 31536 4616
rect 34152 4607 34204 4616
rect 34152 4573 34161 4607
rect 34161 4573 34195 4607
rect 34195 4573 34204 4607
rect 34152 4564 34204 4573
rect 34612 4564 34664 4616
rect 34704 4564 34756 4616
rect 37832 4641 37841 4675
rect 37841 4641 37875 4675
rect 37875 4641 37884 4675
rect 37832 4632 37884 4641
rect 23204 4428 23256 4480
rect 23480 4428 23532 4480
rect 27160 4428 27212 4480
rect 27712 4428 27764 4480
rect 29644 4428 29696 4480
rect 32220 4471 32272 4480
rect 32220 4437 32229 4471
rect 32229 4437 32263 4471
rect 32263 4437 32272 4471
rect 32220 4428 32272 4437
rect 32680 4471 32732 4480
rect 32680 4437 32689 4471
rect 32689 4437 32723 4471
rect 32723 4437 32732 4471
rect 32680 4428 32732 4437
rect 34428 4428 34480 4480
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 19984 4224 20036 4276
rect 21456 4156 21508 4208
rect 21732 4156 21784 4208
rect 20628 4088 20680 4140
rect 21640 4131 21692 4140
rect 21640 4097 21649 4131
rect 21649 4097 21683 4131
rect 21683 4097 21692 4131
rect 21640 4088 21692 4097
rect 22468 4088 22520 4140
rect 24860 4224 24912 4276
rect 25412 4224 25464 4276
rect 26976 4224 27028 4276
rect 27804 4224 27856 4276
rect 28448 4224 28500 4276
rect 28632 4224 28684 4276
rect 29552 4267 29604 4276
rect 29552 4233 29561 4267
rect 29561 4233 29595 4267
rect 29595 4233 29604 4267
rect 29552 4224 29604 4233
rect 30472 4224 30524 4276
rect 33048 4224 33100 4276
rect 34152 4224 34204 4276
rect 34336 4224 34388 4276
rect 34704 4224 34756 4276
rect 35256 4267 35308 4276
rect 35256 4233 35265 4267
rect 35265 4233 35299 4267
rect 35299 4233 35308 4267
rect 35256 4224 35308 4233
rect 26884 4131 26936 4140
rect 26884 4097 26893 4131
rect 26893 4097 26927 4131
rect 26927 4097 26936 4131
rect 26884 4088 26936 4097
rect 27620 4088 27672 4140
rect 27804 4131 27856 4140
rect 27804 4097 27813 4131
rect 27813 4097 27847 4131
rect 27847 4097 27856 4131
rect 27804 4088 27856 4097
rect 33508 4156 33560 4208
rect 31484 4131 31536 4140
rect 31484 4097 31493 4131
rect 31493 4097 31527 4131
rect 31527 4097 31536 4131
rect 31484 4088 31536 4097
rect 32036 4088 32088 4140
rect 15568 4063 15620 4072
rect 15568 4029 15577 4063
rect 15577 4029 15611 4063
rect 15611 4029 15620 4063
rect 15568 4020 15620 4029
rect 17224 4020 17276 4072
rect 17500 4020 17552 4072
rect 19892 4063 19944 4072
rect 19892 4029 19901 4063
rect 19901 4029 19935 4063
rect 19935 4029 19944 4063
rect 19892 4020 19944 4029
rect 31852 4020 31904 4072
rect 34796 4063 34848 4072
rect 34796 4029 34805 4063
rect 34805 4029 34839 4063
rect 34839 4029 34848 4063
rect 34796 4020 34848 4029
rect 36084 4063 36136 4072
rect 36084 4029 36093 4063
rect 36093 4029 36127 4063
rect 36127 4029 36136 4063
rect 36084 4020 36136 4029
rect 36360 4020 36412 4072
rect 17960 3952 18012 4004
rect 19248 3952 19300 4004
rect 21456 3952 21508 4004
rect 25320 3952 25372 4004
rect 16396 3927 16448 3936
rect 16396 3893 16405 3927
rect 16405 3893 16439 3927
rect 16439 3893 16448 3927
rect 16396 3884 16448 3893
rect 18604 3884 18656 3936
rect 22192 3884 22244 3936
rect 25688 3884 25740 3936
rect 28724 3952 28776 4004
rect 31024 3952 31076 4004
rect 31208 3952 31260 4004
rect 36820 4020 36872 4072
rect 37832 4020 37884 4072
rect 31576 3884 31628 3936
rect 32404 3884 32456 3936
rect 33508 3884 33560 3936
rect 37004 3952 37056 4004
rect 34612 3884 34664 3936
rect 36544 3927 36596 3936
rect 36544 3893 36553 3927
rect 36553 3893 36587 3927
rect 36587 3893 36596 3927
rect 36544 3884 36596 3893
rect 36820 3884 36872 3936
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 18604 3680 18656 3732
rect 19064 3723 19116 3732
rect 19064 3689 19073 3723
rect 19073 3689 19107 3723
rect 19107 3689 19116 3723
rect 19064 3680 19116 3689
rect 16120 3612 16172 3664
rect 14648 3476 14700 3528
rect 17500 3612 17552 3664
rect 18052 3612 18104 3664
rect 25320 3680 25372 3732
rect 28448 3680 28500 3732
rect 28632 3723 28684 3732
rect 28632 3689 28641 3723
rect 28641 3689 28675 3723
rect 28675 3689 28684 3723
rect 28632 3680 28684 3689
rect 28724 3680 28776 3732
rect 31208 3680 31260 3732
rect 21916 3612 21968 3664
rect 22928 3612 22980 3664
rect 25780 3655 25832 3664
rect 22560 3587 22612 3596
rect 17684 3476 17736 3528
rect 17960 3476 18012 3528
rect 20352 3519 20404 3528
rect 16856 3451 16908 3460
rect 16856 3417 16865 3451
rect 16865 3417 16899 3451
rect 16899 3417 16908 3451
rect 16856 3408 16908 3417
rect 20352 3485 20361 3519
rect 20361 3485 20395 3519
rect 20395 3485 20404 3519
rect 22560 3553 22569 3587
rect 22569 3553 22603 3587
rect 22603 3553 22612 3587
rect 22560 3544 22612 3553
rect 25780 3621 25789 3655
rect 25789 3621 25823 3655
rect 25823 3621 25832 3655
rect 25780 3612 25832 3621
rect 25872 3655 25924 3664
rect 25872 3621 25881 3655
rect 25881 3621 25915 3655
rect 25915 3621 25924 3655
rect 27160 3655 27212 3664
rect 25872 3612 25924 3621
rect 27160 3621 27169 3655
rect 27169 3621 27203 3655
rect 27203 3621 27212 3655
rect 27160 3612 27212 3621
rect 29644 3612 29696 3664
rect 36820 3680 36872 3732
rect 37004 3680 37056 3732
rect 37464 3723 37516 3732
rect 31852 3612 31904 3664
rect 20352 3476 20404 3485
rect 19432 3408 19484 3460
rect 24308 3519 24360 3528
rect 24308 3485 24317 3519
rect 24317 3485 24351 3519
rect 24351 3485 24360 3519
rect 24308 3476 24360 3485
rect 26884 3587 26936 3596
rect 26884 3553 26893 3587
rect 26893 3553 26927 3587
rect 26927 3553 26936 3587
rect 26884 3544 26936 3553
rect 28448 3544 28500 3596
rect 29092 3544 29144 3596
rect 29368 3544 29420 3596
rect 31576 3476 31628 3528
rect 31852 3476 31904 3528
rect 33140 3612 33192 3664
rect 34152 3655 34204 3664
rect 34152 3621 34161 3655
rect 34161 3621 34195 3655
rect 34195 3621 34204 3655
rect 34152 3612 34204 3621
rect 35992 3655 36044 3664
rect 35992 3621 36001 3655
rect 36001 3621 36035 3655
rect 36035 3621 36044 3655
rect 35992 3612 36044 3621
rect 36452 3612 36504 3664
rect 33600 3476 33652 3528
rect 34704 3544 34756 3596
rect 37464 3689 37473 3723
rect 37473 3689 37507 3723
rect 37507 3689 37516 3723
rect 37464 3680 37516 3689
rect 37924 3723 37976 3732
rect 37924 3689 37933 3723
rect 37933 3689 37967 3723
rect 37967 3689 37976 3723
rect 37924 3680 37976 3689
rect 17224 3340 17276 3392
rect 22008 3340 22060 3392
rect 23388 3340 23440 3392
rect 24768 3340 24820 3392
rect 28724 3408 28776 3460
rect 28816 3408 28868 3460
rect 28540 3340 28592 3392
rect 29184 3340 29236 3392
rect 32312 3340 32364 3392
rect 32680 3383 32732 3392
rect 32680 3349 32689 3383
rect 32689 3349 32723 3383
rect 32723 3349 32732 3383
rect 32680 3340 32732 3349
rect 32956 3340 33008 3392
rect 34060 3340 34112 3392
rect 35440 3340 35492 3392
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 17684 3179 17736 3188
rect 16488 3068 16540 3120
rect 17684 3145 17693 3179
rect 17693 3145 17727 3179
rect 17727 3145 17736 3179
rect 17684 3136 17736 3145
rect 21548 3136 21600 3188
rect 22836 3136 22888 3188
rect 27712 3136 27764 3188
rect 23020 3068 23072 3120
rect 14648 2975 14700 2984
rect 14648 2941 14657 2975
rect 14657 2941 14691 2975
rect 14691 2941 14700 2975
rect 14648 2932 14700 2941
rect 15200 2864 15252 2916
rect 16488 2864 16540 2916
rect 21364 3000 21416 3052
rect 21732 3000 21784 3052
rect 24032 3043 24084 3052
rect 24032 3009 24041 3043
rect 24041 3009 24075 3043
rect 24075 3009 24084 3043
rect 24032 3000 24084 3009
rect 25136 3043 25188 3052
rect 25136 3009 25145 3043
rect 25145 3009 25179 3043
rect 25179 3009 25188 3043
rect 25136 3000 25188 3009
rect 27528 3000 27580 3052
rect 19432 2975 19484 2984
rect 19432 2941 19441 2975
rect 19441 2941 19475 2975
rect 19475 2941 19484 2975
rect 19892 2975 19944 2984
rect 19432 2932 19484 2941
rect 19892 2941 19901 2975
rect 19901 2941 19935 2975
rect 19935 2941 19944 2975
rect 19892 2932 19944 2941
rect 29184 3136 29236 3188
rect 30656 3136 30708 3188
rect 31300 3136 31352 3188
rect 31576 3136 31628 3188
rect 32680 3136 32732 3188
rect 33048 3179 33100 3188
rect 33048 3145 33057 3179
rect 33057 3145 33091 3179
rect 33091 3145 33100 3179
rect 33048 3136 33100 3145
rect 34152 3136 34204 3188
rect 27988 3068 28040 3120
rect 18696 2864 18748 2916
rect 19064 2864 19116 2916
rect 22008 2864 22060 2916
rect 28540 2932 28592 2984
rect 28908 2932 28960 2984
rect 31300 2975 31352 2984
rect 23940 2796 23992 2848
rect 30656 2864 30708 2916
rect 31300 2941 31309 2975
rect 31309 2941 31343 2975
rect 31343 2941 31352 2975
rect 31300 2932 31352 2941
rect 31484 3000 31536 3052
rect 32956 2932 33008 2984
rect 32772 2864 32824 2916
rect 30288 2796 30340 2848
rect 31484 2796 31536 2848
rect 32956 2796 33008 2848
rect 35348 3000 35400 3052
rect 34796 2975 34848 2984
rect 34796 2941 34805 2975
rect 34805 2941 34839 2975
rect 34839 2941 34848 2975
rect 35440 2975 35492 2984
rect 34796 2932 34848 2941
rect 35440 2941 35449 2975
rect 35449 2941 35483 2975
rect 35483 2941 35492 2975
rect 35440 2932 35492 2941
rect 35532 2975 35584 2984
rect 35532 2941 35541 2975
rect 35541 2941 35575 2975
rect 35575 2941 35584 2975
rect 36452 3043 36504 3052
rect 36452 3009 36461 3043
rect 36461 3009 36495 3043
rect 36495 3009 36504 3043
rect 36452 3000 36504 3009
rect 35532 2932 35584 2941
rect 33140 2864 33192 2916
rect 34520 2907 34572 2916
rect 34520 2873 34529 2907
rect 34529 2873 34563 2907
rect 34563 2873 34572 2907
rect 34520 2864 34572 2873
rect 36728 2975 36780 2984
rect 36728 2941 36737 2975
rect 36737 2941 36771 2975
rect 36771 2941 36780 2975
rect 36728 2932 36780 2941
rect 34612 2796 34664 2848
rect 34704 2796 34756 2848
rect 36452 2796 36504 2848
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 16028 2635 16080 2644
rect 16028 2601 16037 2635
rect 16037 2601 16071 2635
rect 16071 2601 16080 2635
rect 16028 2592 16080 2601
rect 16488 2635 16540 2644
rect 16488 2601 16497 2635
rect 16497 2601 16531 2635
rect 16531 2601 16540 2635
rect 16488 2592 16540 2601
rect 16580 2592 16632 2644
rect 18236 2592 18288 2644
rect 19340 2635 19392 2644
rect 19340 2601 19349 2635
rect 19349 2601 19383 2635
rect 19383 2601 19392 2635
rect 19340 2592 19392 2601
rect 17408 2524 17460 2576
rect 17868 2567 17920 2576
rect 17868 2533 17877 2567
rect 17877 2533 17911 2567
rect 17911 2533 17920 2567
rect 17868 2524 17920 2533
rect 21180 2592 21232 2644
rect 24124 2592 24176 2644
rect 24952 2592 25004 2644
rect 26700 2592 26752 2644
rect 27528 2592 27580 2644
rect 31760 2592 31812 2644
rect 20996 2524 21048 2576
rect 23480 2524 23532 2576
rect 28816 2524 28868 2576
rect 29920 2524 29972 2576
rect 34152 2592 34204 2644
rect 35532 2592 35584 2644
rect 32956 2524 33008 2576
rect 34336 2524 34388 2576
rect 36452 2567 36504 2576
rect 36452 2533 36461 2567
rect 36461 2533 36495 2567
rect 36495 2533 36504 2567
rect 36452 2524 36504 2533
rect 13176 2499 13228 2508
rect 13176 2465 13185 2499
rect 13185 2465 13219 2499
rect 13219 2465 13228 2499
rect 13176 2456 13228 2465
rect 16580 2388 16632 2440
rect 14924 2363 14976 2372
rect 14924 2329 14933 2363
rect 14933 2329 14967 2363
rect 14967 2329 14976 2363
rect 14924 2320 14976 2329
rect 13360 2295 13412 2304
rect 13360 2261 13369 2295
rect 13369 2261 13403 2295
rect 13403 2261 13412 2295
rect 13360 2252 13412 2261
rect 14004 2295 14056 2304
rect 14004 2261 14013 2295
rect 14013 2261 14047 2295
rect 14047 2261 14056 2295
rect 14004 2252 14056 2261
rect 19892 2456 19944 2508
rect 22560 2456 22612 2508
rect 24308 2456 24360 2508
rect 27804 2456 27856 2508
rect 17500 2388 17552 2440
rect 20536 2431 20588 2440
rect 20536 2397 20545 2431
rect 20545 2397 20579 2431
rect 20579 2397 20588 2431
rect 20536 2388 20588 2397
rect 24860 2388 24912 2440
rect 25688 2388 25740 2440
rect 33600 2499 33652 2508
rect 33600 2465 33609 2499
rect 33609 2465 33643 2499
rect 33643 2465 33652 2499
rect 33600 2456 33652 2465
rect 36912 2456 36964 2508
rect 37832 2499 37884 2508
rect 37832 2465 37841 2499
rect 37841 2465 37875 2499
rect 37875 2465 37884 2499
rect 37832 2456 37884 2465
rect 32864 2388 32916 2440
rect 33508 2320 33560 2372
rect 35256 2320 35308 2372
rect 25228 2252 25280 2304
rect 37004 2295 37056 2304
rect 37004 2261 37013 2295
rect 37013 2261 37047 2295
rect 37047 2261 37056 2295
rect 37004 2252 37056 2261
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
rect 13360 2048 13412 2100
rect 20536 2048 20588 2100
rect 22008 2048 22060 2100
rect 37004 2048 37056 2100
rect 14004 1980 14056 2032
rect 20996 1980 21048 2032
rect 24308 1980 24360 2032
rect 13176 1912 13228 1964
rect 24952 1912 25004 1964
rect 29092 1980 29144 2032
rect 34336 1980 34388 2032
rect 31116 1912 31168 1964
<< metal2 >>
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 38106 20088 38162 20097
rect 38106 20023 38162 20032
rect 38120 19922 38148 20023
rect 38108 19916 38160 19922
rect 38108 19858 38160 19864
rect 35256 19712 35308 19718
rect 35256 19654 35308 19660
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 35268 13530 35296 19654
rect 35256 13524 35308 13530
rect 35256 13466 35308 13472
rect 33048 13456 33100 13462
rect 33048 13398 33100 13404
rect 32220 13184 32272 13190
rect 32220 13126 32272 13132
rect 32956 13184 33008 13190
rect 32956 13126 33008 13132
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 31852 12844 31904 12850
rect 31852 12786 31904 12792
rect 30656 12776 30708 12782
rect 30656 12718 30708 12724
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 30668 12306 30696 12718
rect 30656 12300 30708 12306
rect 30656 12242 30708 12248
rect 31864 12238 31892 12786
rect 32232 12306 32260 13126
rect 32968 12782 32996 13126
rect 32956 12776 33008 12782
rect 32956 12718 33008 12724
rect 33060 12646 33088 13398
rect 33416 13320 33468 13326
rect 33416 13262 33468 13268
rect 33428 12986 33456 13262
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 33416 12980 33468 12986
rect 33416 12922 33468 12928
rect 35268 12714 35296 13466
rect 35256 12708 35308 12714
rect 35256 12650 35308 12656
rect 32680 12640 32732 12646
rect 32680 12582 32732 12588
rect 33048 12640 33100 12646
rect 33048 12582 33100 12588
rect 32220 12300 32272 12306
rect 32220 12242 32272 12248
rect 31852 12232 31904 12238
rect 31852 12174 31904 12180
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 27712 11212 27764 11218
rect 27712 11154 27764 11160
rect 23664 11076 23716 11082
rect 23664 11018 23716 11024
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 22836 10124 22888 10130
rect 22836 10066 22888 10072
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 4988 9444 5040 9450
rect 4988 9386 5040 9392
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 5000 800 5028 9386
rect 16028 7268 16080 7274
rect 16028 7210 16080 7216
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 14660 2990 14688 3470
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 15212 2922 15240 4966
rect 15580 4078 15608 5714
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15200 2916 15252 2922
rect 15200 2858 15252 2864
rect 16040 2650 16068 7210
rect 16132 3670 16160 9658
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 20720 9036 20772 9042
rect 20720 8978 20772 8984
rect 20444 8560 20496 8566
rect 20444 8502 20496 8508
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 18972 8084 19024 8090
rect 18972 8026 19024 8032
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 16408 3369 16436 3878
rect 16394 3360 16450 3369
rect 16394 3295 16450 3304
rect 16500 3126 16528 6666
rect 17500 5568 17552 5574
rect 17500 5510 17552 5516
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 16854 3496 16910 3505
rect 16854 3431 16856 3440
rect 16908 3431 16910 3440
rect 16856 3402 16908 3408
rect 17236 3398 17264 4014
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 16488 3120 16540 3126
rect 16488 3062 16540 3068
rect 16488 2916 16540 2922
rect 16488 2858 16540 2864
rect 16500 2650 16528 2858
rect 17328 2774 17356 5306
rect 17512 5234 17540 5510
rect 17500 5228 17552 5234
rect 17500 5170 17552 5176
rect 17512 4758 17540 5170
rect 17500 4752 17552 4758
rect 17500 4694 17552 4700
rect 17512 4078 17540 4694
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 17512 3670 17540 4014
rect 17500 3664 17552 3670
rect 17500 3606 17552 3612
rect 17328 2746 17448 2774
rect 16028 2644 16080 2650
rect 16028 2586 16080 2592
rect 16488 2644 16540 2650
rect 16488 2586 16540 2592
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 13176 2508 13228 2514
rect 13176 2450 13228 2456
rect 13188 1970 13216 2450
rect 16592 2446 16620 2586
rect 17420 2582 17448 2746
rect 17408 2576 17460 2582
rect 17408 2518 17460 2524
rect 17512 2446 17540 3606
rect 17604 3233 17632 4558
rect 17684 3528 17736 3534
rect 17684 3470 17736 3476
rect 17590 3224 17646 3233
rect 17696 3194 17724 3470
rect 17590 3159 17646 3168
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17880 2582 17908 7346
rect 18248 5778 18276 7686
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18236 5772 18288 5778
rect 18236 5714 18288 5720
rect 18052 4480 18104 4486
rect 18052 4422 18104 4428
rect 17960 4004 18012 4010
rect 17960 3946 18012 3952
rect 17972 3534 18000 3946
rect 18064 3670 18092 4422
rect 18052 3664 18104 3670
rect 18052 3606 18104 3612
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 18248 2650 18276 5714
rect 18604 3936 18656 3942
rect 18604 3878 18656 3884
rect 18616 3738 18644 3878
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 18708 2922 18736 6054
rect 18892 5574 18920 6190
rect 18880 5568 18932 5574
rect 18880 5510 18932 5516
rect 18892 4826 18920 5510
rect 18880 4820 18932 4826
rect 18880 4762 18932 4768
rect 18984 3618 19012 8026
rect 19432 8016 19484 8022
rect 19432 7958 19484 7964
rect 19064 6180 19116 6186
rect 19064 6122 19116 6128
rect 19076 3738 19104 6122
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19352 4826 19380 5306
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19156 4480 19208 4486
rect 19156 4422 19208 4428
rect 19064 3732 19116 3738
rect 19064 3674 19116 3680
rect 19168 3641 19196 4422
rect 19246 4040 19302 4049
rect 19246 3975 19248 3984
rect 19300 3975 19302 3984
rect 19248 3946 19300 3952
rect 19444 3754 19472 7958
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 19904 6254 19932 6734
rect 19892 6248 19944 6254
rect 19892 6190 19944 6196
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 19904 5710 19932 6190
rect 20088 5846 20116 7142
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20076 5840 20128 5846
rect 20076 5782 20128 5788
rect 20272 5778 20300 6394
rect 20260 5772 20312 5778
rect 20260 5714 20312 5720
rect 19892 5704 19944 5710
rect 19892 5646 19944 5652
rect 19904 5234 19932 5646
rect 19892 5228 19944 5234
rect 19892 5170 19944 5176
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 19904 4078 19932 5170
rect 20456 5098 20484 8502
rect 20732 7426 20760 8978
rect 20640 7398 20760 7426
rect 20640 7342 20668 7398
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20444 5092 20496 5098
rect 20444 5034 20496 5040
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19996 4282 20024 4966
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 19892 4072 19944 4078
rect 19892 4014 19944 4020
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 19260 3726 19472 3754
rect 19154 3632 19210 3641
rect 18984 3590 19104 3618
rect 19076 2922 19104 3590
rect 19154 3567 19210 3576
rect 19260 3346 19288 3726
rect 20364 3534 20392 4558
rect 20640 4146 20668 5646
rect 21180 5568 21232 5574
rect 21180 5510 21232 5516
rect 21192 5234 21220 5510
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 19432 3460 19484 3466
rect 19432 3402 19484 3408
rect 19260 3318 19380 3346
rect 18696 2916 18748 2922
rect 18696 2858 18748 2864
rect 19064 2916 19116 2922
rect 19064 2858 19116 2864
rect 19352 2650 19380 3318
rect 19444 2990 19472 3402
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19892 2984 19944 2990
rect 19892 2926 19944 2932
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 18236 2644 18288 2650
rect 18236 2586 18288 2592
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 17868 2576 17920 2582
rect 17868 2518 17920 2524
rect 19904 2514 19932 2926
rect 21284 2774 21312 9318
rect 22848 9178 22876 10066
rect 23112 9648 23164 9654
rect 23112 9590 23164 9596
rect 22928 9512 22980 9518
rect 22928 9454 22980 9460
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 22008 8356 22060 8362
rect 22008 8298 22060 8304
rect 21548 7948 21600 7954
rect 21548 7890 21600 7896
rect 21560 7750 21588 7890
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 21456 7472 21508 7478
rect 21456 7414 21508 7420
rect 21364 7336 21416 7342
rect 21468 7290 21496 7414
rect 21416 7284 21496 7290
rect 21364 7278 21496 7284
rect 21376 7262 21496 7278
rect 21364 5908 21416 5914
rect 21364 5850 21416 5856
rect 21376 3058 21404 5850
rect 21468 4826 21496 7262
rect 21824 7200 21876 7206
rect 21824 7142 21876 7148
rect 21640 5636 21692 5642
rect 21640 5578 21692 5584
rect 21548 5024 21600 5030
rect 21548 4966 21600 4972
rect 21456 4820 21508 4826
rect 21456 4762 21508 4768
rect 21468 4214 21496 4762
rect 21456 4208 21508 4214
rect 21456 4150 21508 4156
rect 21456 4004 21508 4010
rect 21456 3946 21508 3952
rect 21468 3913 21496 3946
rect 21454 3904 21510 3913
rect 21454 3839 21510 3848
rect 21560 3194 21588 4966
rect 21652 4146 21680 5578
rect 21730 5400 21786 5409
rect 21730 5335 21732 5344
rect 21784 5335 21786 5344
rect 21732 5306 21784 5312
rect 21732 4208 21784 4214
rect 21732 4150 21784 4156
rect 21640 4140 21692 4146
rect 21640 4082 21692 4088
rect 21548 3188 21600 3194
rect 21548 3130 21600 3136
rect 21744 3058 21772 4150
rect 21836 3777 21864 7142
rect 21822 3768 21878 3777
rect 21822 3703 21878 3712
rect 21928 3670 21956 7686
rect 21916 3664 21968 3670
rect 21916 3606 21968 3612
rect 22020 3398 22048 8298
rect 22388 7886 22416 9114
rect 22940 8430 22968 9454
rect 22928 8424 22980 8430
rect 22928 8366 22980 8372
rect 22376 7880 22428 7886
rect 22376 7822 22428 7828
rect 22468 7812 22520 7818
rect 22468 7754 22520 7760
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 22112 6322 22140 7278
rect 22374 6760 22430 6769
rect 22374 6695 22430 6704
rect 22192 6656 22244 6662
rect 22192 6598 22244 6604
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 22100 6180 22152 6186
rect 22100 6122 22152 6128
rect 22112 4622 22140 6122
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 22204 3942 22232 6598
rect 22388 6458 22416 6695
rect 22376 6452 22428 6458
rect 22376 6394 22428 6400
rect 22480 5166 22508 7754
rect 22940 7342 22968 8366
rect 23020 8288 23072 8294
rect 23020 8230 23072 8236
rect 23032 8022 23060 8230
rect 23020 8016 23072 8022
rect 23020 7958 23072 7964
rect 22928 7336 22980 7342
rect 22928 7278 22980 7284
rect 23020 7336 23072 7342
rect 23020 7278 23072 7284
rect 22560 6792 22612 6798
rect 22560 6734 22612 6740
rect 22572 6322 22600 6734
rect 22928 6656 22980 6662
rect 22928 6598 22980 6604
rect 22560 6316 22612 6322
rect 22560 6258 22612 6264
rect 22572 5778 22600 6258
rect 22560 5772 22612 5778
rect 22560 5714 22612 5720
rect 22834 5264 22890 5273
rect 22834 5199 22836 5208
rect 22888 5199 22890 5208
rect 22836 5170 22888 5176
rect 22468 5160 22520 5166
rect 22468 5102 22520 5108
rect 22834 5128 22890 5137
rect 22480 4146 22508 5102
rect 22834 5063 22836 5072
rect 22888 5063 22890 5072
rect 22836 5034 22888 5040
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 22836 4616 22888 4622
rect 22836 4558 22888 4564
rect 22468 4140 22520 4146
rect 22468 4082 22520 4088
rect 22192 3936 22244 3942
rect 22192 3878 22244 3884
rect 22572 3602 22600 4558
rect 22560 3596 22612 3602
rect 22560 3538 22612 3544
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 21364 3052 21416 3058
rect 21364 2994 21416 3000
rect 21732 3052 21784 3058
rect 21732 2994 21784 3000
rect 22008 2916 22060 2922
rect 22008 2858 22060 2864
rect 21192 2746 21312 2774
rect 21192 2650 21220 2746
rect 21180 2644 21232 2650
rect 21180 2586 21232 2592
rect 20996 2576 21048 2582
rect 20996 2518 21048 2524
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 16580 2440 16632 2446
rect 16580 2382 16632 2388
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 14924 2372 14976 2378
rect 14924 2314 14976 2320
rect 13360 2304 13412 2310
rect 13360 2246 13412 2252
rect 14004 2304 14056 2310
rect 14004 2246 14056 2252
rect 13372 2106 13400 2246
rect 13360 2100 13412 2106
rect 13360 2042 13412 2048
rect 14016 2038 14044 2246
rect 14004 2032 14056 2038
rect 14004 1974 14056 1980
rect 13176 1964 13228 1970
rect 13176 1906 13228 1912
rect 14936 800 14964 2314
rect 20548 2106 20576 2382
rect 20536 2100 20588 2106
rect 20536 2042 20588 2048
rect 21008 2038 21036 2518
rect 22020 2106 22048 2858
rect 22572 2514 22600 3538
rect 22848 3194 22876 4558
rect 22940 3670 22968 6598
rect 22928 3664 22980 3670
rect 22928 3606 22980 3612
rect 22836 3188 22888 3194
rect 22836 3130 22888 3136
rect 23032 3126 23060 7278
rect 23124 6934 23152 9590
rect 23676 9042 23704 11018
rect 24124 10736 24176 10742
rect 24124 10678 24176 10684
rect 23664 9036 23716 9042
rect 23664 8978 23716 8984
rect 23676 8922 23704 8978
rect 23584 8894 23704 8922
rect 23848 8968 23900 8974
rect 23848 8910 23900 8916
rect 23480 8288 23532 8294
rect 23480 8230 23532 8236
rect 23112 6928 23164 6934
rect 23112 6870 23164 6876
rect 23388 5704 23440 5710
rect 23388 5646 23440 5652
rect 23112 5364 23164 5370
rect 23112 5306 23164 5312
rect 23124 4758 23152 5306
rect 23112 4752 23164 4758
rect 23112 4694 23164 4700
rect 23204 4616 23256 4622
rect 23204 4558 23256 4564
rect 23216 4486 23244 4558
rect 23204 4480 23256 4486
rect 23204 4422 23256 4428
rect 23400 3398 23428 5646
rect 23492 4622 23520 8230
rect 23584 7750 23612 8894
rect 23664 8832 23716 8838
rect 23664 8774 23716 8780
rect 23572 7744 23624 7750
rect 23572 7686 23624 7692
rect 23676 5098 23704 8774
rect 23860 8430 23888 8910
rect 23848 8424 23900 8430
rect 23848 8366 23900 8372
rect 23940 7336 23992 7342
rect 23940 7278 23992 7284
rect 23664 5092 23716 5098
rect 23664 5034 23716 5040
rect 23480 4616 23532 4622
rect 23480 4558 23532 4564
rect 23480 4480 23532 4486
rect 23480 4422 23532 4428
rect 23388 3392 23440 3398
rect 23388 3334 23440 3340
rect 23020 3120 23072 3126
rect 23020 3062 23072 3068
rect 23492 2582 23520 4422
rect 23952 2854 23980 7278
rect 24136 5846 24164 10678
rect 27252 10668 27304 10674
rect 27252 10610 27304 10616
rect 25872 10124 25924 10130
rect 25872 10066 25924 10072
rect 24952 9988 25004 9994
rect 24952 9930 25004 9936
rect 24308 9920 24360 9926
rect 24308 9862 24360 9868
rect 24320 8566 24348 9862
rect 24676 9512 24728 9518
rect 24676 9454 24728 9460
rect 24308 8560 24360 8566
rect 24308 8502 24360 8508
rect 24320 7954 24348 8502
rect 24400 8356 24452 8362
rect 24400 8298 24452 8304
rect 24308 7948 24360 7954
rect 24308 7890 24360 7896
rect 24320 7410 24348 7890
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 24216 6860 24268 6866
rect 24216 6802 24268 6808
rect 24228 6769 24256 6802
rect 24412 6798 24440 8298
rect 24688 8294 24716 9454
rect 24768 8832 24820 8838
rect 24768 8774 24820 8780
rect 24676 8288 24728 8294
rect 24676 8230 24728 8236
rect 24584 7404 24636 7410
rect 24584 7346 24636 7352
rect 24400 6792 24452 6798
rect 24214 6760 24270 6769
rect 24400 6734 24452 6740
rect 24214 6695 24270 6704
rect 24492 6384 24544 6390
rect 24596 6372 24624 7346
rect 24544 6344 24624 6372
rect 24492 6326 24544 6332
rect 24596 6254 24624 6344
rect 24584 6248 24636 6254
rect 24584 6190 24636 6196
rect 24124 5840 24176 5846
rect 24124 5782 24176 5788
rect 24308 5636 24360 5642
rect 24308 5578 24360 5584
rect 24032 5568 24084 5574
rect 24032 5510 24084 5516
rect 24044 3058 24072 5510
rect 24124 5092 24176 5098
rect 24124 5034 24176 5040
rect 24032 3052 24084 3058
rect 24032 2994 24084 3000
rect 23940 2848 23992 2854
rect 23940 2790 23992 2796
rect 24136 2650 24164 5034
rect 24320 3534 24348 5578
rect 24308 3528 24360 3534
rect 24308 3470 24360 3476
rect 24780 3398 24808 8774
rect 24860 7268 24912 7274
rect 24860 7210 24912 7216
rect 24872 5914 24900 7210
rect 24964 6390 24992 9930
rect 25780 9920 25832 9926
rect 25780 9862 25832 9868
rect 25792 9722 25820 9862
rect 25780 9716 25832 9722
rect 25780 9658 25832 9664
rect 25884 9518 25912 10066
rect 26700 9988 26752 9994
rect 26700 9930 26752 9936
rect 26332 9920 26384 9926
rect 26332 9862 26384 9868
rect 25872 9512 25924 9518
rect 25872 9454 25924 9460
rect 25412 9376 25464 9382
rect 25412 9318 25464 9324
rect 25424 9110 25452 9318
rect 25412 9104 25464 9110
rect 25412 9046 25464 9052
rect 26240 9104 26292 9110
rect 26240 9046 26292 9052
rect 25044 8832 25096 8838
rect 25044 8774 25096 8780
rect 24952 6384 25004 6390
rect 24952 6326 25004 6332
rect 24952 6180 25004 6186
rect 24952 6122 25004 6128
rect 24860 5908 24912 5914
rect 24860 5850 24912 5856
rect 24860 4276 24912 4282
rect 24860 4218 24912 4224
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24124 2644 24176 2650
rect 24124 2586 24176 2592
rect 23480 2576 23532 2582
rect 23480 2518 23532 2524
rect 22560 2508 22612 2514
rect 22560 2450 22612 2456
rect 24308 2508 24360 2514
rect 24308 2450 24360 2456
rect 22008 2100 22060 2106
rect 22008 2042 22060 2048
rect 24320 2038 24348 2450
rect 24872 2446 24900 4218
rect 24964 2650 24992 6122
rect 25056 5137 25084 8774
rect 25228 8288 25280 8294
rect 25228 8230 25280 8236
rect 25240 6730 25268 8230
rect 25504 7880 25556 7886
rect 25504 7822 25556 7828
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 25228 6724 25280 6730
rect 25228 6666 25280 6672
rect 25240 6361 25268 6666
rect 25226 6352 25282 6361
rect 25226 6287 25282 6296
rect 25136 5296 25188 5302
rect 25136 5238 25188 5244
rect 25148 5166 25176 5238
rect 25136 5160 25188 5166
rect 25042 5128 25098 5137
rect 25136 5102 25188 5108
rect 25042 5063 25098 5072
rect 25148 4690 25176 5102
rect 25136 4684 25188 4690
rect 25136 4626 25188 4632
rect 25148 3058 25176 4626
rect 25136 3052 25188 3058
rect 25136 2994 25188 3000
rect 24952 2644 25004 2650
rect 24952 2586 25004 2592
rect 24860 2440 24912 2446
rect 24860 2382 24912 2388
rect 25240 2310 25268 6287
rect 25424 5710 25452 7482
rect 25516 6458 25544 7822
rect 26252 7546 26280 9046
rect 26240 7540 26292 7546
rect 26240 7482 26292 7488
rect 25780 7200 25832 7206
rect 25780 7142 25832 7148
rect 25504 6452 25556 6458
rect 25504 6394 25556 6400
rect 25412 5704 25464 5710
rect 25412 5646 25464 5652
rect 25412 5092 25464 5098
rect 25412 5034 25464 5040
rect 25424 4282 25452 5034
rect 25504 5024 25556 5030
rect 25504 4966 25556 4972
rect 25516 4758 25544 4966
rect 25504 4752 25556 4758
rect 25504 4694 25556 4700
rect 25412 4276 25464 4282
rect 25412 4218 25464 4224
rect 25320 4004 25372 4010
rect 25320 3946 25372 3952
rect 25332 3738 25360 3946
rect 25688 3936 25740 3942
rect 25688 3878 25740 3884
rect 25320 3732 25372 3738
rect 25320 3674 25372 3680
rect 25700 2446 25728 3878
rect 25792 3670 25820 7142
rect 25872 5704 25924 5710
rect 25872 5646 25924 5652
rect 25884 3670 25912 5646
rect 26344 5273 26372 9862
rect 26424 7200 26476 7206
rect 26424 7142 26476 7148
rect 26436 6934 26464 7142
rect 26424 6928 26476 6934
rect 26424 6870 26476 6876
rect 26330 5264 26386 5273
rect 26330 5199 26386 5208
rect 25780 3664 25832 3670
rect 25780 3606 25832 3612
rect 25872 3664 25924 3670
rect 25872 3606 25924 3612
rect 26712 2650 26740 9930
rect 27264 9382 27292 10610
rect 27724 10130 27752 11154
rect 31864 11150 31892 12174
rect 32692 11286 32720 12582
rect 33060 12374 33088 12582
rect 33048 12368 33100 12374
rect 33048 12310 33100 12316
rect 33048 12096 33100 12102
rect 33048 12038 33100 12044
rect 32680 11280 32732 11286
rect 32680 11222 32732 11228
rect 33060 11218 33088 12038
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 33048 11212 33100 11218
rect 33048 11154 33100 11160
rect 31852 11144 31904 11150
rect 31852 11086 31904 11092
rect 31392 11076 31444 11082
rect 31392 11018 31444 11024
rect 27896 10600 27948 10606
rect 27896 10542 27948 10548
rect 30840 10600 30892 10606
rect 30840 10542 30892 10548
rect 27804 10464 27856 10470
rect 27804 10406 27856 10412
rect 27712 10124 27764 10130
rect 27712 10066 27764 10072
rect 27528 9580 27580 9586
rect 27528 9522 27580 9528
rect 27436 9444 27488 9450
rect 27436 9386 27488 9392
rect 27252 9376 27304 9382
rect 27252 9318 27304 9324
rect 27264 8906 27292 9318
rect 27252 8900 27304 8906
rect 27252 8842 27304 8848
rect 26976 7744 27028 7750
rect 26976 7686 27028 7692
rect 26988 4282 27016 7686
rect 27158 5808 27214 5817
rect 27158 5743 27160 5752
rect 27212 5743 27214 5752
rect 27160 5714 27212 5720
rect 27160 4480 27212 4486
rect 27160 4422 27212 4428
rect 26976 4276 27028 4282
rect 26976 4218 27028 4224
rect 26884 4140 26936 4146
rect 26884 4082 26936 4088
rect 26896 3602 26924 4082
rect 27172 3670 27200 4422
rect 27264 4321 27292 8842
rect 27344 6792 27396 6798
rect 27344 6734 27396 6740
rect 27356 6662 27384 6734
rect 27344 6656 27396 6662
rect 27344 6598 27396 6604
rect 27356 6066 27384 6598
rect 27448 6186 27476 9386
rect 27436 6180 27488 6186
rect 27436 6122 27488 6128
rect 27434 6080 27490 6089
rect 27356 6038 27434 6066
rect 27434 6015 27490 6024
rect 27448 5642 27476 6015
rect 27436 5636 27488 5642
rect 27436 5578 27488 5584
rect 27436 5228 27488 5234
rect 27436 5170 27488 5176
rect 27448 4758 27476 5170
rect 27540 5098 27568 9522
rect 27620 9512 27672 9518
rect 27620 9454 27672 9460
rect 27632 9042 27660 9454
rect 27620 9036 27672 9042
rect 27620 8978 27672 8984
rect 27632 6662 27660 8978
rect 27724 8634 27752 10066
rect 27816 8974 27844 10406
rect 27908 8974 27936 10542
rect 28908 10192 28960 10198
rect 28908 10134 28960 10140
rect 28080 10056 28132 10062
rect 28080 9998 28132 10004
rect 28092 9042 28120 9998
rect 28724 9648 28776 9654
rect 28724 9590 28776 9596
rect 28540 9376 28592 9382
rect 28540 9318 28592 9324
rect 28080 9036 28132 9042
rect 28080 8978 28132 8984
rect 27804 8968 27856 8974
rect 27804 8910 27856 8916
rect 27896 8968 27948 8974
rect 27896 8910 27948 8916
rect 27712 8628 27764 8634
rect 27712 8570 27764 8576
rect 27816 8378 27844 8910
rect 28092 8838 28120 8978
rect 28080 8832 28132 8838
rect 28080 8774 28132 8780
rect 28172 8832 28224 8838
rect 28172 8774 28224 8780
rect 27724 8350 27844 8378
rect 27896 8356 27948 8362
rect 27724 7886 27752 8350
rect 27896 8298 27948 8304
rect 27804 8288 27856 8294
rect 27804 8230 27856 8236
rect 27816 8022 27844 8230
rect 27804 8016 27856 8022
rect 27804 7958 27856 7964
rect 27712 7880 27764 7886
rect 27712 7822 27764 7828
rect 27724 6662 27752 7822
rect 27908 7750 27936 8298
rect 28092 7886 28120 8774
rect 28080 7880 28132 7886
rect 28080 7822 28132 7828
rect 27896 7744 27948 7750
rect 27896 7686 27948 7692
rect 27896 7200 27948 7206
rect 27896 7142 27948 7148
rect 27804 6792 27856 6798
rect 27804 6734 27856 6740
rect 27620 6656 27672 6662
rect 27620 6598 27672 6604
rect 27712 6656 27764 6662
rect 27712 6598 27764 6604
rect 27620 6384 27672 6390
rect 27620 6326 27672 6332
rect 27632 6100 27660 6326
rect 27724 6254 27752 6598
rect 27712 6248 27764 6254
rect 27712 6190 27764 6196
rect 27816 6100 27844 6734
rect 27632 6072 27844 6100
rect 27804 5568 27856 5574
rect 27804 5510 27856 5516
rect 27528 5092 27580 5098
rect 27528 5034 27580 5040
rect 27712 5024 27764 5030
rect 27712 4966 27764 4972
rect 27724 4758 27752 4966
rect 27436 4752 27488 4758
rect 27436 4694 27488 4700
rect 27712 4752 27764 4758
rect 27712 4694 27764 4700
rect 27436 4616 27488 4622
rect 27488 4564 27660 4570
rect 27436 4558 27660 4564
rect 27448 4542 27660 4558
rect 27250 4312 27306 4321
rect 27250 4247 27306 4256
rect 27632 4146 27660 4542
rect 27712 4480 27764 4486
rect 27712 4422 27764 4428
rect 27620 4140 27672 4146
rect 27620 4082 27672 4088
rect 27160 3664 27212 3670
rect 27160 3606 27212 3612
rect 26884 3596 26936 3602
rect 26884 3538 26936 3544
rect 27724 3194 27752 4422
rect 27816 4282 27844 5510
rect 27908 5409 27936 7142
rect 28184 7002 28212 8774
rect 28446 8528 28502 8537
rect 28446 8463 28502 8472
rect 28172 6996 28224 7002
rect 28172 6938 28224 6944
rect 28460 6610 28488 8463
rect 28552 7274 28580 9318
rect 28632 8016 28684 8022
rect 28632 7958 28684 7964
rect 28644 7410 28672 7958
rect 28632 7404 28684 7410
rect 28632 7346 28684 7352
rect 28540 7268 28592 7274
rect 28540 7210 28592 7216
rect 28644 6882 28672 7346
rect 28552 6866 28672 6882
rect 28540 6860 28672 6866
rect 28592 6854 28672 6860
rect 28540 6802 28592 6808
rect 28368 6582 28488 6610
rect 28078 6352 28134 6361
rect 28078 6287 28080 6296
rect 28132 6287 28134 6296
rect 28080 6258 28132 6264
rect 28080 6180 28132 6186
rect 28080 6122 28132 6128
rect 28092 5710 28120 6122
rect 28080 5704 28132 5710
rect 28080 5646 28132 5652
rect 27988 5568 28040 5574
rect 27988 5510 28040 5516
rect 27894 5400 27950 5409
rect 27894 5335 27950 5344
rect 27804 4276 27856 4282
rect 27804 4218 27856 4224
rect 27804 4140 27856 4146
rect 28000 4128 28028 5510
rect 28368 4758 28396 6582
rect 28448 5704 28500 5710
rect 28448 5646 28500 5652
rect 28356 4752 28408 4758
rect 28356 4694 28408 4700
rect 28460 4282 28488 5646
rect 28448 4276 28500 4282
rect 28448 4218 28500 4224
rect 27856 4100 28028 4128
rect 27804 4082 27856 4088
rect 27712 3188 27764 3194
rect 27712 3130 27764 3136
rect 28000 3126 28028 4100
rect 28448 3732 28500 3738
rect 28448 3674 28500 3680
rect 28460 3602 28488 3674
rect 28448 3596 28500 3602
rect 28448 3538 28500 3544
rect 28552 3398 28580 6802
rect 28632 4276 28684 4282
rect 28632 4218 28684 4224
rect 28644 3738 28672 4218
rect 28736 4010 28764 9590
rect 28920 9518 28948 10134
rect 30852 10130 30880 10542
rect 31024 10532 31076 10538
rect 31024 10474 31076 10480
rect 30840 10124 30892 10130
rect 30840 10066 30892 10072
rect 29920 10056 29972 10062
rect 29920 9998 29972 10004
rect 29092 9920 29144 9926
rect 29092 9862 29144 9868
rect 29104 9518 29132 9862
rect 29932 9518 29960 9998
rect 30656 9920 30708 9926
rect 30656 9862 30708 9868
rect 28908 9512 28960 9518
rect 28908 9454 28960 9460
rect 29092 9512 29144 9518
rect 29092 9454 29144 9460
rect 29920 9512 29972 9518
rect 29920 9454 29972 9460
rect 28920 9042 28948 9454
rect 29104 9042 29132 9454
rect 30472 9444 30524 9450
rect 30472 9386 30524 9392
rect 29184 9376 29236 9382
rect 29184 9318 29236 9324
rect 28908 9036 28960 9042
rect 28908 8978 28960 8984
rect 29092 9036 29144 9042
rect 29092 8978 29144 8984
rect 28920 8945 28948 8978
rect 28906 8936 28962 8945
rect 28906 8871 28962 8880
rect 28908 8832 28960 8838
rect 28908 8774 28960 8780
rect 28816 8492 28868 8498
rect 28816 8434 28868 8440
rect 28828 6202 28856 8434
rect 28920 6934 28948 8774
rect 29196 8650 29224 9318
rect 30288 9104 30340 9110
rect 30288 9046 30340 9052
rect 30196 9036 30248 9042
rect 30196 8978 30248 8984
rect 30104 8968 30156 8974
rect 30104 8910 30156 8916
rect 29104 8622 29224 8650
rect 30116 8634 30144 8910
rect 30104 8628 30156 8634
rect 28908 6928 28960 6934
rect 28908 6870 28960 6876
rect 28828 6174 28948 6202
rect 28816 6112 28868 6118
rect 28816 6054 28868 6060
rect 28828 5710 28856 6054
rect 28816 5704 28868 5710
rect 28816 5646 28868 5652
rect 28814 5264 28870 5273
rect 28814 5199 28816 5208
rect 28868 5199 28870 5208
rect 28816 5170 28868 5176
rect 28920 5114 28948 6174
rect 28998 5808 29054 5817
rect 28998 5743 29000 5752
rect 29052 5743 29054 5752
rect 29000 5714 29052 5720
rect 28920 5098 29040 5114
rect 28920 5092 29052 5098
rect 28920 5086 29000 5092
rect 29000 5034 29052 5040
rect 28724 4004 28776 4010
rect 28724 3946 28776 3952
rect 28632 3732 28684 3738
rect 28632 3674 28684 3680
rect 28724 3732 28776 3738
rect 28724 3674 28776 3680
rect 28736 3466 28764 3674
rect 29104 3602 29132 8622
rect 30104 8570 30156 8576
rect 29552 8560 29604 8566
rect 29550 8528 29552 8537
rect 29604 8528 29606 8537
rect 29184 8492 29236 8498
rect 29550 8463 29606 8472
rect 29184 8434 29236 8440
rect 29196 4622 29224 8434
rect 29552 8424 29604 8430
rect 29552 8366 29604 8372
rect 29564 7342 29592 8366
rect 30208 7886 30236 8978
rect 30196 7880 30248 7886
rect 30196 7822 30248 7828
rect 29920 7472 29972 7478
rect 29920 7414 29972 7420
rect 29552 7336 29604 7342
rect 29550 7304 29552 7313
rect 29604 7304 29606 7313
rect 29550 7239 29606 7248
rect 29564 6866 29592 7239
rect 29826 7032 29882 7041
rect 29826 6967 29882 6976
rect 29552 6860 29604 6866
rect 29552 6802 29604 6808
rect 29276 6656 29328 6662
rect 29276 6598 29328 6604
rect 29184 4616 29236 4622
rect 29184 4558 29236 4564
rect 29092 3596 29144 3602
rect 29092 3538 29144 3544
rect 28724 3460 28776 3466
rect 28724 3402 28776 3408
rect 28816 3460 28868 3466
rect 28816 3402 28868 3408
rect 28540 3392 28592 3398
rect 28540 3334 28592 3340
rect 27988 3120 28040 3126
rect 27988 3062 28040 3068
rect 27528 3052 27580 3058
rect 27528 2994 27580 3000
rect 27540 2650 27568 2994
rect 28000 2774 28028 3062
rect 28552 2990 28580 3334
rect 28540 2984 28592 2990
rect 28540 2926 28592 2932
rect 27816 2746 28028 2774
rect 26700 2644 26752 2650
rect 26700 2586 26752 2592
rect 27528 2644 27580 2650
rect 27528 2586 27580 2592
rect 27816 2514 27844 2746
rect 28828 2582 28856 3402
rect 29184 3392 29236 3398
rect 29184 3334 29236 3340
rect 29196 3194 29224 3334
rect 29184 3188 29236 3194
rect 29184 3130 29236 3136
rect 28906 3088 28962 3097
rect 28906 3023 28962 3032
rect 28920 2990 28948 3023
rect 28908 2984 28960 2990
rect 28908 2926 28960 2932
rect 29288 2774 29316 6598
rect 29458 6352 29514 6361
rect 29458 6287 29460 6296
rect 29512 6287 29514 6296
rect 29460 6258 29512 6264
rect 29368 5568 29420 5574
rect 29368 5510 29420 5516
rect 29380 3602 29408 5510
rect 29564 5234 29592 6802
rect 29840 5574 29868 6967
rect 29828 5568 29880 5574
rect 29828 5510 29880 5516
rect 29644 5296 29696 5302
rect 29644 5238 29696 5244
rect 29734 5264 29790 5273
rect 29552 5228 29604 5234
rect 29552 5170 29604 5176
rect 29656 4570 29684 5238
rect 29734 5199 29736 5208
rect 29788 5199 29790 5208
rect 29736 5170 29788 5176
rect 29564 4542 29684 4570
rect 29564 4282 29592 4542
rect 29644 4480 29696 4486
rect 29644 4422 29696 4428
rect 29552 4276 29604 4282
rect 29552 4218 29604 4224
rect 29656 3670 29684 4422
rect 29644 3664 29696 3670
rect 29644 3606 29696 3612
rect 29368 3596 29420 3602
rect 29368 3538 29420 3544
rect 29104 2746 29316 2774
rect 28816 2576 28868 2582
rect 28816 2518 28868 2524
rect 27804 2508 27856 2514
rect 27804 2450 27856 2456
rect 25688 2440 25740 2446
rect 25688 2382 25740 2388
rect 25228 2304 25280 2310
rect 25228 2246 25280 2252
rect 29104 2038 29132 2746
rect 29932 2582 29960 7414
rect 30208 7410 30236 7822
rect 30196 7404 30248 7410
rect 30196 7346 30248 7352
rect 30196 7200 30248 7206
rect 30196 7142 30248 7148
rect 30012 6996 30064 7002
rect 30012 6938 30064 6944
rect 30024 5642 30052 6938
rect 30208 6934 30236 7142
rect 30196 6928 30248 6934
rect 30196 6870 30248 6876
rect 30196 6180 30248 6186
rect 30196 6122 30248 6128
rect 30104 6112 30156 6118
rect 30104 6054 30156 6060
rect 30116 5914 30144 6054
rect 30104 5908 30156 5914
rect 30104 5850 30156 5856
rect 30208 5642 30236 6122
rect 30300 5914 30328 9046
rect 30484 8906 30512 9386
rect 30668 9042 30696 9862
rect 30656 9036 30708 9042
rect 30656 8978 30708 8984
rect 30654 8936 30710 8945
rect 30472 8900 30524 8906
rect 30852 8906 30880 10066
rect 30654 8871 30710 8880
rect 30840 8900 30892 8906
rect 30472 8842 30524 8848
rect 30380 8832 30432 8838
rect 30380 8774 30432 8780
rect 30288 5908 30340 5914
rect 30288 5850 30340 5856
rect 30392 5778 30420 8774
rect 30668 7954 30696 8871
rect 30840 8842 30892 8848
rect 30656 7948 30708 7954
rect 30656 7890 30708 7896
rect 30668 7206 30696 7890
rect 30840 7812 30892 7818
rect 30840 7754 30892 7760
rect 30932 7812 30984 7818
rect 30932 7754 30984 7760
rect 30748 7540 30800 7546
rect 30748 7482 30800 7488
rect 30656 7200 30708 7206
rect 30656 7142 30708 7148
rect 30760 6746 30788 7482
rect 30852 7342 30880 7754
rect 30944 7478 30972 7754
rect 30932 7472 30984 7478
rect 30932 7414 30984 7420
rect 30840 7336 30892 7342
rect 30840 7278 30892 7284
rect 30932 7336 30984 7342
rect 30932 7278 30984 7284
rect 30944 7206 30972 7278
rect 30932 7200 30984 7206
rect 30932 7142 30984 7148
rect 30576 6718 30788 6746
rect 30472 6384 30524 6390
rect 30472 6326 30524 6332
rect 30380 5772 30432 5778
rect 30380 5714 30432 5720
rect 30012 5636 30064 5642
rect 30012 5578 30064 5584
rect 30196 5636 30248 5642
rect 30196 5578 30248 5584
rect 30024 4758 30052 5578
rect 30380 5092 30432 5098
rect 30380 5034 30432 5040
rect 30012 4752 30064 4758
rect 30012 4694 30064 4700
rect 30392 4690 30420 5034
rect 30380 4684 30432 4690
rect 30380 4626 30432 4632
rect 30286 4448 30342 4457
rect 30286 4383 30342 4392
rect 30300 2854 30328 4383
rect 30484 4282 30512 6326
rect 30576 5098 30604 6718
rect 30656 6656 30708 6662
rect 30656 6598 30708 6604
rect 30564 5092 30616 5098
rect 30564 5034 30616 5040
rect 30472 4276 30524 4282
rect 30472 4218 30524 4224
rect 30668 3194 30696 6598
rect 30748 6316 30800 6322
rect 30748 6258 30800 6264
rect 30760 4758 30788 6258
rect 31036 6186 31064 10474
rect 31208 10056 31260 10062
rect 31208 9998 31260 10004
rect 31220 8634 31248 9998
rect 31208 8628 31260 8634
rect 31208 8570 31260 8576
rect 31116 7744 31168 7750
rect 31116 7686 31168 7692
rect 31024 6180 31076 6186
rect 31024 6122 31076 6128
rect 31022 5264 31078 5273
rect 31022 5199 31078 5208
rect 30748 4752 30800 4758
rect 30748 4694 30800 4700
rect 31036 4010 31064 5199
rect 31024 4004 31076 4010
rect 31024 3946 31076 3952
rect 30656 3188 30708 3194
rect 30656 3130 30708 3136
rect 30668 2922 30696 3130
rect 30656 2916 30708 2922
rect 30656 2858 30708 2864
rect 30288 2848 30340 2854
rect 30288 2790 30340 2796
rect 29920 2576 29972 2582
rect 29920 2518 29972 2524
rect 20996 2032 21048 2038
rect 20996 1974 21048 1980
rect 24308 2032 24360 2038
rect 24308 1974 24360 1980
rect 29092 2032 29144 2038
rect 29092 1974 29144 1980
rect 31128 1970 31156 7686
rect 31220 5817 31248 8570
rect 31404 8430 31432 11018
rect 31864 10266 31892 11086
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 31852 10260 31904 10266
rect 31852 10202 31904 10208
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 32036 9580 32088 9586
rect 32036 9522 32088 9528
rect 31668 9512 31720 9518
rect 31668 9454 31720 9460
rect 31484 8968 31536 8974
rect 31484 8910 31536 8916
rect 31392 8424 31444 8430
rect 31392 8366 31444 8372
rect 31496 8294 31524 8910
rect 31680 8430 31708 9454
rect 31668 8424 31720 8430
rect 31668 8366 31720 8372
rect 31484 8288 31536 8294
rect 31484 8230 31536 8236
rect 31576 7880 31628 7886
rect 31576 7822 31628 7828
rect 31392 7336 31444 7342
rect 31392 7278 31444 7284
rect 31300 7200 31352 7206
rect 31300 7142 31352 7148
rect 31206 5808 31262 5817
rect 31206 5743 31262 5752
rect 31312 5098 31340 7142
rect 31300 5092 31352 5098
rect 31300 5034 31352 5040
rect 31208 4004 31260 4010
rect 31208 3946 31260 3952
rect 31220 3738 31248 3946
rect 31208 3732 31260 3738
rect 31208 3674 31260 3680
rect 31300 3188 31352 3194
rect 31300 3130 31352 3136
rect 31312 2990 31340 3130
rect 31404 3040 31432 7278
rect 31588 7002 31616 7822
rect 31680 7041 31708 8366
rect 32048 7954 32076 9522
rect 37832 9036 37884 9042
rect 37832 8978 37884 8984
rect 35440 8832 35492 8838
rect 35440 8774 35492 8780
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 32496 8016 32548 8022
rect 32496 7958 32548 7964
rect 32036 7948 32088 7954
rect 32036 7890 32088 7896
rect 31852 7744 31904 7750
rect 31852 7686 31904 7692
rect 31666 7032 31722 7041
rect 31576 6996 31628 7002
rect 31666 6967 31722 6976
rect 31576 6938 31628 6944
rect 31668 6928 31720 6934
rect 31496 6876 31668 6882
rect 31496 6870 31720 6876
rect 31496 6854 31708 6870
rect 31496 6798 31524 6854
rect 31864 6798 31892 7686
rect 31944 7200 31996 7206
rect 31944 7142 31996 7148
rect 31484 6792 31536 6798
rect 31484 6734 31536 6740
rect 31576 6792 31628 6798
rect 31576 6734 31628 6740
rect 31852 6792 31904 6798
rect 31852 6734 31904 6740
rect 31484 6180 31536 6186
rect 31484 6122 31536 6128
rect 31496 4729 31524 6122
rect 31588 5914 31616 6734
rect 31760 6656 31812 6662
rect 31760 6598 31812 6604
rect 31666 6216 31722 6225
rect 31666 6151 31722 6160
rect 31576 5908 31628 5914
rect 31576 5850 31628 5856
rect 31482 4720 31538 4729
rect 31482 4655 31538 4664
rect 31484 4616 31536 4622
rect 31484 4558 31536 4564
rect 31496 4146 31524 4558
rect 31574 4176 31630 4185
rect 31484 4140 31536 4146
rect 31574 4111 31630 4120
rect 31484 4082 31536 4088
rect 31588 3942 31616 4111
rect 31576 3936 31628 3942
rect 31576 3878 31628 3884
rect 31576 3528 31628 3534
rect 31680 3516 31708 6151
rect 31772 4593 31800 6598
rect 31852 6452 31904 6458
rect 31852 6394 31904 6400
rect 31864 6322 31892 6394
rect 31852 6316 31904 6322
rect 31852 6258 31904 6264
rect 31850 5944 31906 5953
rect 31850 5879 31906 5888
rect 31864 5846 31892 5879
rect 31852 5840 31904 5846
rect 31852 5782 31904 5788
rect 31758 4584 31814 4593
rect 31758 4519 31814 4528
rect 31956 4185 31984 7142
rect 32048 7002 32076 7890
rect 32402 7304 32458 7313
rect 32402 7239 32458 7248
rect 32310 7032 32366 7041
rect 32036 6996 32088 7002
rect 32310 6967 32366 6976
rect 32036 6938 32088 6944
rect 32324 6866 32352 6967
rect 32312 6860 32364 6866
rect 32312 6802 32364 6808
rect 32416 6798 32444 7239
rect 32404 6792 32456 6798
rect 32404 6734 32456 6740
rect 32220 6452 32272 6458
rect 32220 6394 32272 6400
rect 32312 6452 32364 6458
rect 32312 6394 32364 6400
rect 32036 6384 32088 6390
rect 32036 6326 32088 6332
rect 32048 6225 32076 6326
rect 32128 6248 32180 6254
rect 32034 6216 32090 6225
rect 32128 6190 32180 6196
rect 32034 6151 32090 6160
rect 32140 6089 32168 6190
rect 32126 6080 32182 6089
rect 32126 6015 32182 6024
rect 32232 5710 32260 6394
rect 32220 5704 32272 5710
rect 32220 5646 32272 5652
rect 32232 5166 32260 5646
rect 32220 5160 32272 5166
rect 32220 5102 32272 5108
rect 32220 5024 32272 5030
rect 32220 4966 32272 4972
rect 32232 4486 32260 4966
rect 32220 4480 32272 4486
rect 32220 4422 32272 4428
rect 32034 4312 32090 4321
rect 32034 4247 32090 4256
rect 31942 4176 31998 4185
rect 32048 4146 32076 4247
rect 31942 4111 31998 4120
rect 32036 4140 32088 4146
rect 32036 4082 32088 4088
rect 31852 4072 31904 4078
rect 31852 4014 31904 4020
rect 31864 3670 31892 4014
rect 31852 3664 31904 3670
rect 31852 3606 31904 3612
rect 31628 3488 31708 3516
rect 31852 3528 31904 3534
rect 31576 3470 31628 3476
rect 31852 3470 31904 3476
rect 31576 3188 31628 3194
rect 31576 3130 31628 3136
rect 31588 3097 31616 3130
rect 31574 3088 31630 3097
rect 31484 3052 31536 3058
rect 31404 3012 31484 3040
rect 31574 3023 31630 3032
rect 31484 2994 31536 3000
rect 31300 2984 31352 2990
rect 31300 2926 31352 2932
rect 31484 2848 31536 2854
rect 31482 2816 31484 2825
rect 31536 2816 31538 2825
rect 31482 2751 31538 2760
rect 31864 2666 31892 3470
rect 32324 3398 32352 6394
rect 32508 5098 32536 7958
rect 32692 6866 32720 8434
rect 33140 8288 33192 8294
rect 33140 8230 33192 8236
rect 33152 7954 33180 8230
rect 33140 7948 33192 7954
rect 33140 7890 33192 7896
rect 34612 7948 34664 7954
rect 34612 7890 34664 7896
rect 33152 7342 33180 7890
rect 33140 7336 33192 7342
rect 33140 7278 33192 7284
rect 33692 7336 33744 7342
rect 33692 7278 33744 7284
rect 32956 7268 33008 7274
rect 32956 7210 33008 7216
rect 32680 6860 32732 6866
rect 32680 6802 32732 6808
rect 32772 6656 32824 6662
rect 32772 6598 32824 6604
rect 32784 5846 32812 6598
rect 32862 6352 32918 6361
rect 32862 6287 32918 6296
rect 32772 5840 32824 5846
rect 32772 5782 32824 5788
rect 32876 5778 32904 6287
rect 32968 6254 32996 7210
rect 33048 6860 33100 6866
rect 33048 6802 33100 6808
rect 33416 6860 33468 6866
rect 33416 6802 33468 6808
rect 32956 6248 33008 6254
rect 32956 6190 33008 6196
rect 32968 5778 32996 6190
rect 33060 5914 33088 6802
rect 33140 6724 33192 6730
rect 33140 6666 33192 6672
rect 33048 5908 33100 5914
rect 33048 5850 33100 5856
rect 32864 5772 32916 5778
rect 32864 5714 32916 5720
rect 32956 5772 33008 5778
rect 32956 5714 33008 5720
rect 32772 5568 32824 5574
rect 32772 5510 32824 5516
rect 32496 5092 32548 5098
rect 32496 5034 32548 5040
rect 32678 4720 32734 4729
rect 32678 4655 32734 4664
rect 32692 4486 32720 4655
rect 32680 4480 32732 4486
rect 32680 4422 32732 4428
rect 32404 3936 32456 3942
rect 32404 3878 32456 3884
rect 32312 3392 32364 3398
rect 32312 3334 32364 3340
rect 32416 3233 32444 3878
rect 32680 3392 32732 3398
rect 32680 3334 32732 3340
rect 32402 3224 32458 3233
rect 32692 3194 32720 3334
rect 32402 3159 32458 3168
rect 32680 3188 32732 3194
rect 32680 3130 32732 3136
rect 32784 2922 32812 5510
rect 33048 5296 33100 5302
rect 33152 5250 33180 6666
rect 33428 5574 33456 6802
rect 33324 5568 33376 5574
rect 33324 5510 33376 5516
rect 33416 5568 33468 5574
rect 33416 5510 33468 5516
rect 33100 5244 33180 5250
rect 33048 5238 33180 5244
rect 33060 5222 33180 5238
rect 33048 5160 33100 5166
rect 33046 5128 33048 5137
rect 33100 5128 33102 5137
rect 33046 5063 33102 5072
rect 32864 4752 32916 4758
rect 32864 4694 32916 4700
rect 32772 2916 32824 2922
rect 32772 2858 32824 2864
rect 31772 2650 31892 2666
rect 31760 2644 31892 2650
rect 31812 2638 31892 2644
rect 31760 2586 31812 2592
rect 32876 2446 32904 4694
rect 33048 4276 33100 4282
rect 33048 4218 33100 4224
rect 32956 3392 33008 3398
rect 32956 3334 33008 3340
rect 32968 2990 32996 3334
rect 33060 3194 33088 4218
rect 33336 4049 33364 5510
rect 33508 4208 33560 4214
rect 33508 4150 33560 4156
rect 33322 4040 33378 4049
rect 33322 3975 33378 3984
rect 33520 3942 33548 4150
rect 33508 3936 33560 3942
rect 33508 3878 33560 3884
rect 33138 3768 33194 3777
rect 33138 3703 33194 3712
rect 33506 3768 33562 3777
rect 33506 3703 33562 3712
rect 33152 3670 33180 3703
rect 33140 3664 33192 3670
rect 33140 3606 33192 3612
rect 33138 3360 33194 3369
rect 33138 3295 33194 3304
rect 33048 3188 33100 3194
rect 33048 3130 33100 3136
rect 32956 2984 33008 2990
rect 32956 2926 33008 2932
rect 33152 2922 33180 3295
rect 33140 2916 33192 2922
rect 33140 2858 33192 2864
rect 32956 2848 33008 2854
rect 32956 2790 33008 2796
rect 32968 2582 32996 2790
rect 32956 2576 33008 2582
rect 32956 2518 33008 2524
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 33520 2378 33548 3703
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 33612 2514 33640 3470
rect 33704 2825 33732 7278
rect 34152 7268 34204 7274
rect 34152 7210 34204 7216
rect 34060 7200 34112 7206
rect 34060 7142 34112 7148
rect 33876 6248 33928 6254
rect 33876 6190 33928 6196
rect 33888 5846 33916 6190
rect 33876 5840 33928 5846
rect 33876 5782 33928 5788
rect 33784 5092 33836 5098
rect 33784 5034 33836 5040
rect 33796 4457 33824 5034
rect 33782 4448 33838 4457
rect 33782 4383 33838 4392
rect 34072 3398 34100 7142
rect 34164 6866 34192 7210
rect 34624 6866 34652 7890
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 34704 6996 34756 7002
rect 34704 6938 34756 6944
rect 34152 6860 34204 6866
rect 34152 6802 34204 6808
rect 34612 6860 34664 6866
rect 34612 6802 34664 6808
rect 34164 4706 34192 6802
rect 34612 6656 34664 6662
rect 34612 6598 34664 6604
rect 34336 6316 34388 6322
rect 34336 6258 34388 6264
rect 34348 5030 34376 6258
rect 34624 5137 34652 6598
rect 34716 6322 34744 6938
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 34704 6316 34756 6322
rect 34704 6258 34756 6264
rect 35348 6248 35400 6254
rect 35348 6190 35400 6196
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 34610 5128 34666 5137
rect 34610 5063 34666 5072
rect 34244 5024 34296 5030
rect 34244 4966 34296 4972
rect 34336 5024 34388 5030
rect 34336 4966 34388 4972
rect 34256 4842 34284 4966
rect 34256 4814 34560 4842
rect 34164 4678 34284 4706
rect 34532 4690 34560 4814
rect 34152 4616 34204 4622
rect 34152 4558 34204 4564
rect 34164 4282 34192 4558
rect 34152 4276 34204 4282
rect 34256 4264 34284 4678
rect 34520 4684 34572 4690
rect 34520 4626 34572 4632
rect 34624 4622 34652 5063
rect 35256 4752 35308 4758
rect 35256 4694 35308 4700
rect 34612 4616 34664 4622
rect 34612 4558 34664 4564
rect 34704 4616 34756 4622
rect 34704 4558 34756 4564
rect 34428 4480 34480 4486
rect 34428 4422 34480 4428
rect 34336 4276 34388 4282
rect 34256 4236 34336 4264
rect 34152 4218 34204 4224
rect 34336 4218 34388 4224
rect 34440 3777 34468 4422
rect 34624 4060 34652 4558
rect 34716 4282 34744 4558
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 35268 4282 35296 4694
rect 35360 4690 35388 6190
rect 35452 5166 35480 8774
rect 35716 8356 35768 8362
rect 35716 8298 35768 8304
rect 35532 6316 35584 6322
rect 35532 6258 35584 6264
rect 35544 5166 35572 6258
rect 35728 5914 35756 8298
rect 36544 8084 36596 8090
rect 36544 8026 36596 8032
rect 35808 6860 35860 6866
rect 35808 6802 35860 6808
rect 35716 5908 35768 5914
rect 35716 5850 35768 5856
rect 35716 5364 35768 5370
rect 35716 5306 35768 5312
rect 35728 5273 35756 5306
rect 35714 5264 35770 5273
rect 35714 5199 35770 5208
rect 35440 5160 35492 5166
rect 35440 5102 35492 5108
rect 35532 5160 35584 5166
rect 35532 5102 35584 5108
rect 35452 4690 35480 5102
rect 35820 4826 35848 6802
rect 35900 6792 35952 6798
rect 35900 6734 35952 6740
rect 35912 5778 35940 6734
rect 36084 6180 36136 6186
rect 36084 6122 36136 6128
rect 35900 5772 35952 5778
rect 35900 5714 35952 5720
rect 35912 5098 35940 5714
rect 35992 5296 36044 5302
rect 35992 5238 36044 5244
rect 35900 5092 35952 5098
rect 35900 5034 35952 5040
rect 35808 4820 35860 4826
rect 35808 4762 35860 4768
rect 35348 4684 35400 4690
rect 35348 4626 35400 4632
rect 35440 4684 35492 4690
rect 35440 4626 35492 4632
rect 34704 4276 34756 4282
rect 34704 4218 34756 4224
rect 35256 4276 35308 4282
rect 35256 4218 35308 4224
rect 34796 4072 34848 4078
rect 34624 4032 34796 4060
rect 34612 3936 34664 3942
rect 34612 3878 34664 3884
rect 34426 3768 34482 3777
rect 34426 3703 34482 3712
rect 34152 3664 34204 3670
rect 34150 3632 34152 3641
rect 34204 3632 34206 3641
rect 34150 3567 34206 3576
rect 34518 3496 34574 3505
rect 34518 3431 34574 3440
rect 34060 3392 34112 3398
rect 34060 3334 34112 3340
rect 34152 3188 34204 3194
rect 34152 3130 34204 3136
rect 33690 2816 33746 2825
rect 33690 2751 33746 2760
rect 34164 2650 34192 3130
rect 34532 2922 34560 3431
rect 34520 2916 34572 2922
rect 34520 2858 34572 2864
rect 34624 2854 34652 3878
rect 34716 3602 34744 4032
rect 34796 4014 34848 4020
rect 34704 3596 34756 3602
rect 34704 3538 34756 3544
rect 34716 2972 34744 3538
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 35360 3058 35388 4626
rect 36004 3670 36032 5238
rect 36096 4078 36124 6122
rect 36452 5568 36504 5574
rect 36452 5510 36504 5516
rect 36360 4684 36412 4690
rect 36360 4626 36412 4632
rect 36372 4078 36400 4626
rect 36084 4072 36136 4078
rect 36084 4014 36136 4020
rect 36360 4072 36412 4078
rect 36360 4014 36412 4020
rect 36464 3670 36492 5510
rect 36556 3942 36584 8026
rect 36912 7404 36964 7410
rect 36912 7346 36964 7352
rect 36728 6112 36780 6118
rect 36728 6054 36780 6060
rect 36544 3936 36596 3942
rect 36544 3878 36596 3884
rect 35992 3664 36044 3670
rect 35992 3606 36044 3612
rect 36452 3664 36504 3670
rect 36452 3606 36504 3612
rect 35440 3392 35492 3398
rect 35440 3334 35492 3340
rect 35348 3052 35400 3058
rect 35348 2994 35400 3000
rect 35452 2990 35480 3334
rect 36452 3052 36504 3058
rect 36452 2994 36504 3000
rect 34796 2984 34848 2990
rect 34716 2944 34796 2972
rect 34796 2926 34848 2932
rect 35440 2984 35492 2990
rect 35440 2926 35492 2932
rect 35532 2984 35584 2990
rect 35532 2926 35584 2932
rect 34612 2848 34664 2854
rect 34704 2848 34756 2854
rect 34612 2790 34664 2796
rect 34702 2816 34704 2825
rect 34756 2816 34758 2825
rect 34702 2751 34758 2760
rect 35544 2650 35572 2926
rect 36464 2854 36492 2994
rect 36740 2990 36768 6054
rect 36820 5704 36872 5710
rect 36820 5646 36872 5652
rect 36832 4690 36860 5646
rect 36820 4684 36872 4690
rect 36820 4626 36872 4632
rect 36832 4078 36860 4626
rect 36820 4072 36872 4078
rect 36820 4014 36872 4020
rect 36820 3936 36872 3942
rect 36820 3878 36872 3884
rect 36832 3738 36860 3878
rect 36820 3732 36872 3738
rect 36820 3674 36872 3680
rect 36728 2984 36780 2990
rect 36728 2926 36780 2932
rect 36452 2848 36504 2854
rect 36452 2790 36504 2796
rect 34152 2644 34204 2650
rect 34152 2586 34204 2592
rect 35532 2644 35584 2650
rect 35532 2586 35584 2592
rect 36464 2582 36492 2790
rect 34336 2576 34388 2582
rect 34336 2518 34388 2524
rect 36452 2576 36504 2582
rect 36452 2518 36504 2524
rect 33600 2508 33652 2514
rect 33600 2450 33652 2456
rect 33508 2372 33560 2378
rect 33508 2314 33560 2320
rect 34348 2038 34376 2518
rect 36924 2514 36952 7346
rect 37844 4690 37872 8978
rect 37832 4684 37884 4690
rect 37832 4626 37884 4632
rect 37462 4584 37518 4593
rect 37462 4519 37518 4528
rect 37004 4004 37056 4010
rect 37004 3946 37056 3952
rect 37016 3738 37044 3946
rect 37476 3738 37504 4519
rect 37832 4072 37884 4078
rect 37832 4014 37884 4020
rect 37004 3732 37056 3738
rect 37004 3674 37056 3680
rect 37464 3732 37516 3738
rect 37464 3674 37516 3680
rect 37844 2514 37872 4014
rect 37922 3904 37978 3913
rect 37922 3839 37978 3848
rect 37936 3738 37964 3839
rect 37924 3732 37976 3738
rect 37924 3674 37976 3680
rect 36912 2508 36964 2514
rect 36912 2450 36964 2456
rect 37832 2508 37884 2514
rect 37832 2450 37884 2456
rect 35256 2372 35308 2378
rect 35256 2314 35308 2320
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 34336 2032 34388 2038
rect 34336 1974 34388 1980
rect 24952 1964 25004 1970
rect 24952 1906 25004 1912
rect 31116 1964 31168 1970
rect 31116 1906 31168 1912
rect 24964 800 24992 1906
rect 35268 1170 35296 2314
rect 37004 2304 37056 2310
rect 37004 2246 37056 2252
rect 37016 2106 37044 2246
rect 37004 2100 37056 2106
rect 37004 2042 37056 2048
rect 34992 1142 35296 1170
rect 34992 800 35020 1142
rect 4986 0 5042 800
rect 14922 0 14978 800
rect 24950 0 25006 800
rect 34978 0 35034 800
<< via2 >>
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 38106 20032 38162 20088
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 16394 3304 16450 3360
rect 16854 3460 16910 3496
rect 16854 3440 16856 3460
rect 16856 3440 16908 3460
rect 16908 3440 16910 3460
rect 17590 3168 17646 3224
rect 19246 4004 19302 4040
rect 19246 3984 19248 4004
rect 19248 3984 19300 4004
rect 19300 3984 19302 4004
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19154 3576 19210 3632
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 21454 3848 21510 3904
rect 21730 5364 21786 5400
rect 21730 5344 21732 5364
rect 21732 5344 21784 5364
rect 21784 5344 21786 5364
rect 21822 3712 21878 3768
rect 22374 6704 22430 6760
rect 22834 5228 22890 5264
rect 22834 5208 22836 5228
rect 22836 5208 22888 5228
rect 22888 5208 22890 5228
rect 22834 5092 22890 5128
rect 22834 5072 22836 5092
rect 22836 5072 22888 5092
rect 22888 5072 22890 5092
rect 24214 6704 24270 6760
rect 25226 6296 25282 6352
rect 25042 5072 25098 5128
rect 26330 5208 26386 5264
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 27158 5772 27214 5808
rect 27158 5752 27160 5772
rect 27160 5752 27212 5772
rect 27212 5752 27214 5772
rect 27434 6024 27490 6080
rect 27250 4256 27306 4312
rect 28446 8472 28502 8528
rect 28078 6316 28134 6352
rect 28078 6296 28080 6316
rect 28080 6296 28132 6316
rect 28132 6296 28134 6316
rect 27894 5344 27950 5400
rect 28906 8880 28962 8936
rect 28814 5228 28870 5264
rect 28814 5208 28816 5228
rect 28816 5208 28868 5228
rect 28868 5208 28870 5228
rect 28998 5772 29054 5808
rect 28998 5752 29000 5772
rect 29000 5752 29052 5772
rect 29052 5752 29054 5772
rect 29550 8508 29552 8528
rect 29552 8508 29604 8528
rect 29604 8508 29606 8528
rect 29550 8472 29606 8508
rect 29550 7284 29552 7304
rect 29552 7284 29604 7304
rect 29604 7284 29606 7304
rect 29550 7248 29606 7284
rect 29826 6976 29882 7032
rect 28906 3032 28962 3088
rect 29458 6316 29514 6352
rect 29458 6296 29460 6316
rect 29460 6296 29512 6316
rect 29512 6296 29514 6316
rect 29734 5228 29790 5264
rect 29734 5208 29736 5228
rect 29736 5208 29788 5228
rect 29788 5208 29790 5228
rect 30654 8880 30710 8936
rect 30286 4392 30342 4448
rect 31022 5208 31078 5264
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 31206 5752 31262 5808
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 31666 6976 31722 7032
rect 31666 6160 31722 6216
rect 31482 4664 31538 4720
rect 31574 4120 31630 4176
rect 31850 5888 31906 5944
rect 31758 4528 31814 4584
rect 32402 7248 32458 7304
rect 32310 6976 32366 7032
rect 32034 6160 32090 6216
rect 32126 6024 32182 6080
rect 32034 4256 32090 4312
rect 31942 4120 31998 4176
rect 31574 3032 31630 3088
rect 31482 2796 31484 2816
rect 31484 2796 31536 2816
rect 31536 2796 31538 2816
rect 31482 2760 31538 2796
rect 32862 6296 32918 6352
rect 32678 4664 32734 4720
rect 32402 3168 32458 3224
rect 33046 5108 33048 5128
rect 33048 5108 33100 5128
rect 33100 5108 33102 5128
rect 33046 5072 33102 5108
rect 33322 3984 33378 4040
rect 33138 3712 33194 3768
rect 33506 3712 33562 3768
rect 33138 3304 33194 3360
rect 33782 4392 33838 4448
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 34610 5072 34666 5128
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 35714 5208 35770 5264
rect 34426 3712 34482 3768
rect 34150 3612 34152 3632
rect 34152 3612 34204 3632
rect 34204 3612 34206 3632
rect 34150 3576 34206 3612
rect 34518 3440 34574 3496
rect 33690 2760 33746 2816
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 34702 2796 34704 2816
rect 34704 2796 34756 2816
rect 34756 2796 34758 2816
rect 34702 2760 34758 2796
rect 37462 4528 37518 4584
rect 37922 3848 37978 3904
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
<< metal3 >>
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 28255 35248 28256
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 27167 35248 27168
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 38101 20090 38167 20093
rect 39200 20090 40000 20120
rect 38101 20088 40000 20090
rect 38101 20032 38106 20088
rect 38162 20032 40000 20088
rect 38101 20030 40000 20032
rect 38101 20027 38167 20030
rect 39200 20000 40000 20030
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 16287 35248 16288
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 13023 35248 13024
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 10847 35248 10848
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 28901 8938 28967 8941
rect 30649 8938 30715 8941
rect 28901 8936 30715 8938
rect 28901 8880 28906 8936
rect 28962 8880 30654 8936
rect 30710 8880 30715 8936
rect 28901 8878 30715 8880
rect 28901 8875 28967 8878
rect 30649 8875 30715 8878
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 28441 8530 28507 8533
rect 29545 8530 29611 8533
rect 28441 8528 29611 8530
rect 28441 8472 28446 8528
rect 28502 8472 29550 8528
rect 29606 8472 29611 8528
rect 28441 8470 29611 8472
rect 28441 8467 28507 8470
rect 29545 8467 29611 8470
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 29545 7306 29611 7309
rect 32397 7306 32463 7309
rect 29545 7304 32463 7306
rect 29545 7248 29550 7304
rect 29606 7248 32402 7304
rect 32458 7248 32463 7304
rect 29545 7246 32463 7248
rect 29545 7243 29611 7246
rect 32397 7243 32463 7246
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 29821 7034 29887 7037
rect 31661 7034 31727 7037
rect 32305 7034 32371 7037
rect 29821 7032 32371 7034
rect 29821 6976 29826 7032
rect 29882 6976 31666 7032
rect 31722 6976 32310 7032
rect 32366 6976 32371 7032
rect 29821 6974 32371 6976
rect 29821 6971 29887 6974
rect 31661 6971 31727 6974
rect 32305 6971 32371 6974
rect 22369 6762 22435 6765
rect 24209 6762 24275 6765
rect 22369 6760 24275 6762
rect 22369 6704 22374 6760
rect 22430 6704 24214 6760
rect 24270 6704 24275 6760
rect 22369 6702 24275 6704
rect 22369 6699 22435 6702
rect 24209 6699 24275 6702
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 6495 35248 6496
rect 25221 6354 25287 6357
rect 28073 6354 28139 6357
rect 25221 6352 28139 6354
rect 25221 6296 25226 6352
rect 25282 6296 28078 6352
rect 28134 6296 28139 6352
rect 25221 6294 28139 6296
rect 25221 6291 25287 6294
rect 28073 6291 28139 6294
rect 29453 6354 29519 6357
rect 32857 6354 32923 6357
rect 29453 6352 32923 6354
rect 29453 6296 29458 6352
rect 29514 6296 32862 6352
rect 32918 6296 32923 6352
rect 29453 6294 32923 6296
rect 29453 6291 29519 6294
rect 32857 6291 32923 6294
rect 31661 6218 31727 6221
rect 32029 6218 32095 6221
rect 31661 6216 32095 6218
rect 31661 6160 31666 6216
rect 31722 6160 32034 6216
rect 32090 6160 32095 6216
rect 31661 6158 32095 6160
rect 31661 6155 31727 6158
rect 32029 6155 32095 6158
rect 27429 6082 27495 6085
rect 32121 6082 32187 6085
rect 27429 6080 32187 6082
rect 27429 6024 27434 6080
rect 27490 6024 32126 6080
rect 32182 6024 32187 6080
rect 27429 6022 32187 6024
rect 27429 6019 27495 6022
rect 32121 6019 32187 6022
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 31845 5946 31911 5949
rect 31710 5944 31911 5946
rect 31710 5888 31850 5944
rect 31906 5888 31911 5944
rect 31710 5886 31911 5888
rect 27153 5810 27219 5813
rect 28993 5810 29059 5813
rect 31201 5810 31267 5813
rect 31710 5810 31770 5886
rect 31845 5883 31911 5886
rect 27153 5808 31770 5810
rect 27153 5752 27158 5808
rect 27214 5752 28998 5808
rect 29054 5752 31206 5808
rect 31262 5752 31770 5808
rect 27153 5750 31770 5752
rect 27153 5747 27219 5750
rect 28993 5747 29059 5750
rect 31201 5747 31267 5750
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 21725 5402 21791 5405
rect 27889 5402 27955 5405
rect 21725 5400 27955 5402
rect 21725 5344 21730 5400
rect 21786 5344 27894 5400
rect 27950 5344 27955 5400
rect 21725 5342 27955 5344
rect 21725 5339 21791 5342
rect 27889 5339 27955 5342
rect 22829 5266 22895 5269
rect 26325 5266 26391 5269
rect 22829 5264 26391 5266
rect 22829 5208 22834 5264
rect 22890 5208 26330 5264
rect 26386 5208 26391 5264
rect 22829 5206 26391 5208
rect 22829 5203 22895 5206
rect 26325 5203 26391 5206
rect 28809 5266 28875 5269
rect 29729 5266 29795 5269
rect 28809 5264 29795 5266
rect 28809 5208 28814 5264
rect 28870 5208 29734 5264
rect 29790 5208 29795 5264
rect 28809 5206 29795 5208
rect 28809 5203 28875 5206
rect 29729 5203 29795 5206
rect 31017 5266 31083 5269
rect 35709 5266 35775 5269
rect 31017 5264 35775 5266
rect 31017 5208 31022 5264
rect 31078 5208 35714 5264
rect 35770 5208 35775 5264
rect 31017 5206 35775 5208
rect 31017 5203 31083 5206
rect 35709 5203 35775 5206
rect 22829 5130 22895 5133
rect 25037 5130 25103 5133
rect 22829 5128 25103 5130
rect 22829 5072 22834 5128
rect 22890 5072 25042 5128
rect 25098 5072 25103 5128
rect 22829 5070 25103 5072
rect 22829 5067 22895 5070
rect 25037 5067 25103 5070
rect 33041 5130 33107 5133
rect 34605 5130 34671 5133
rect 33041 5128 34671 5130
rect 33041 5072 33046 5128
rect 33102 5072 34610 5128
rect 34666 5072 34671 5128
rect 33041 5070 34671 5072
rect 33041 5067 33107 5070
rect 34605 5067 34671 5070
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 31477 4722 31543 4725
rect 32673 4722 32739 4725
rect 31477 4720 32739 4722
rect 31477 4664 31482 4720
rect 31538 4664 32678 4720
rect 32734 4664 32739 4720
rect 31477 4662 32739 4664
rect 31477 4659 31543 4662
rect 32673 4659 32739 4662
rect 31753 4586 31819 4589
rect 37457 4586 37523 4589
rect 31753 4584 37523 4586
rect 31753 4528 31758 4584
rect 31814 4528 37462 4584
rect 37518 4528 37523 4584
rect 31753 4526 37523 4528
rect 31753 4523 31819 4526
rect 37457 4523 37523 4526
rect 30281 4450 30347 4453
rect 33777 4450 33843 4453
rect 30281 4448 33843 4450
rect 30281 4392 30286 4448
rect 30342 4392 33782 4448
rect 33838 4392 33843 4448
rect 30281 4390 33843 4392
rect 30281 4387 30347 4390
rect 33777 4387 33843 4390
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 27245 4314 27311 4317
rect 32029 4314 32095 4317
rect 27245 4312 32095 4314
rect 27245 4256 27250 4312
rect 27306 4256 32034 4312
rect 32090 4256 32095 4312
rect 27245 4254 32095 4256
rect 27245 4251 27311 4254
rect 32029 4251 32095 4254
rect 31569 4178 31635 4181
rect 31937 4178 32003 4181
rect 31569 4176 32003 4178
rect 31569 4120 31574 4176
rect 31630 4120 31942 4176
rect 31998 4120 32003 4176
rect 31569 4118 32003 4120
rect 31569 4115 31635 4118
rect 31937 4115 32003 4118
rect 19241 4042 19307 4045
rect 33317 4042 33383 4045
rect 19241 4040 33383 4042
rect 19241 3984 19246 4040
rect 19302 3984 33322 4040
rect 33378 3984 33383 4040
rect 19241 3982 33383 3984
rect 19241 3979 19307 3982
rect 33317 3979 33383 3982
rect 21449 3906 21515 3909
rect 37917 3906 37983 3909
rect 21449 3904 37983 3906
rect 21449 3848 21454 3904
rect 21510 3848 37922 3904
rect 37978 3848 37983 3904
rect 21449 3846 37983 3848
rect 21449 3843 21515 3846
rect 37917 3843 37983 3846
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 21817 3770 21883 3773
rect 33133 3770 33199 3773
rect 21817 3768 33199 3770
rect 21817 3712 21822 3768
rect 21878 3712 33138 3768
rect 33194 3712 33199 3768
rect 21817 3710 33199 3712
rect 21817 3707 21883 3710
rect 33133 3707 33199 3710
rect 33501 3770 33567 3773
rect 34421 3770 34487 3773
rect 33501 3768 34487 3770
rect 33501 3712 33506 3768
rect 33562 3712 34426 3768
rect 34482 3712 34487 3768
rect 33501 3710 34487 3712
rect 33501 3707 33567 3710
rect 34421 3707 34487 3710
rect 19149 3634 19215 3637
rect 34145 3634 34211 3637
rect 19149 3632 34211 3634
rect 19149 3576 19154 3632
rect 19210 3576 34150 3632
rect 34206 3576 34211 3632
rect 19149 3574 34211 3576
rect 19149 3571 19215 3574
rect 34145 3571 34211 3574
rect 16849 3498 16915 3501
rect 34513 3498 34579 3501
rect 16849 3496 34579 3498
rect 16849 3440 16854 3496
rect 16910 3440 34518 3496
rect 34574 3440 34579 3496
rect 16849 3438 34579 3440
rect 16849 3435 16915 3438
rect 34513 3435 34579 3438
rect 16389 3362 16455 3365
rect 33133 3362 33199 3365
rect 16389 3360 33199 3362
rect 16389 3304 16394 3360
rect 16450 3304 33138 3360
rect 33194 3304 33199 3360
rect 16389 3302 33199 3304
rect 16389 3299 16455 3302
rect 33133 3299 33199 3302
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 17585 3226 17651 3229
rect 32397 3226 32463 3229
rect 17585 3224 32463 3226
rect 17585 3168 17590 3224
rect 17646 3168 32402 3224
rect 32458 3168 32463 3224
rect 17585 3166 32463 3168
rect 17585 3163 17651 3166
rect 32397 3163 32463 3166
rect 28901 3090 28967 3093
rect 31569 3090 31635 3093
rect 28901 3088 31635 3090
rect 28901 3032 28906 3088
rect 28962 3032 31574 3088
rect 31630 3032 31635 3088
rect 28901 3030 31635 3032
rect 28901 3027 28967 3030
rect 31569 3027 31635 3030
rect 31477 2818 31543 2821
rect 33685 2818 33751 2821
rect 34697 2818 34763 2821
rect 31477 2816 34763 2818
rect 31477 2760 31482 2816
rect 31538 2760 33690 2816
rect 33746 2760 34702 2816
rect 34758 2760 34763 2816
rect 31477 2758 34763 2760
rect 31477 2755 31543 2758
rect 33685 2755 33751 2758
rect 34697 2755 34763 2758
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
<< via3 >>
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
<< metal4 >>
rect 4208 37024 4528 37584
rect 19568 37568 19888 37584
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4868 2176 5188 37536
rect 5528 2176 5848 37536
rect 6188 2176 6508 37536
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 4208 2128 4528 2144
rect 19568 2128 19888 2688
rect 20228 2176 20548 37536
rect 20888 2176 21208 37536
rect 21548 2176 21868 37536
rect 34928 37024 35248 37584
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 35588 2176 35908 37536
rect 36248 2176 36568 37536
rect 36908 2176 37228 37536
rect 34928 2128 35248 2144
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1623529830
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1623529830
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1623529830
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1623529830
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_30
timestamp 1623529830
transform 1 0 3864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_42
timestamp 1623529830
transform 1 0 4968 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1623529830
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1623529830
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1623529830
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1623529830
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_59
timestamp 1623529830
transform 1 0 6532 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 5796 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_58
timestamp 1623529830
transform 1 0 6440 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1623529830
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_71
timestamp 1623529830
transform 1 0 7636 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1623529830
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_70
timestamp 1623529830
transform 1 0 7544 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_82
timestamp 1623529830
transform 1 0 8648 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_88
timestamp 1623529830
transform 1 0 9200 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_100
timestamp 1623529830
transform 1 0 10304 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_94
timestamp 1623529830
transform 1 0 9752 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_106 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 10856 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1623529830
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1623529830
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform -1 0 13432 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1623529830
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_117
timestamp 1623529830
transform 1 0 11868 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_129
timestamp 1623529830
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_115
timestamp 1623529830
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_127
timestamp 1623529830
transform 1 0 12788 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_139 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 13892 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1623529830
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_134
timestamp 1623529830
transform 1 0 13432 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _168_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform -1 0 14260 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp 1623529830
transform -1 0 14076 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_143
timestamp 1623529830
transform 1 0 14260 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1623529830
transform 1 0 14536 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform -1 0 15272 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1623529830
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _235_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 14628 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1623529830
transform 1 0 16468 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _136_
timestamp 1623529830
transform -1 0 16100 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1623529830
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1623529830
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_154
timestamp 1623529830
transform 1 0 15272 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1623529830
transform 1 0 16100 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_170
timestamp 1623529830
transform 1 0 16744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_167
timestamp 1623529830
transform 1 0 16468 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_172
timestamp 1623529830
transform 1 0 16928 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _224_
timestamp 1623529830
transform -1 0 19504 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _226_
timestamp 1623529830
transform 1 0 17572 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1623529830
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _202_
timestamp 1623529830
transform 1 0 19872 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _204_
timestamp 1623529830
transform 1 0 20240 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1623529830
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_199
timestamp 1623529830
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_204
timestamp 1623529830
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_200
timestamp 1623529830
transform 1 0 19504 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _200_
timestamp 1623529830
transform 1 0 22908 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _205_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform -1 0 24472 0 1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1623529830
transform 1 0 22448 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1623529830
transform 1 0 22080 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_228
timestamp 1623529830
transform 1 0 22080 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_233
timestamp 1623529830
transform 1 0 22540 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_224
timestamp 1623529830
transform 1 0 21712 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_229
timestamp 1623529830
transform 1 0 22172 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _189_
timestamp 1623529830
transform 1 0 25116 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1623529830
transform 1 0 25116 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_257
timestamp 1623529830
transform 1 0 24748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1623529830
transform 1 0 25208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_254
timestamp 1623529830
transform 1 0 24472 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_260
timestamp 1623529830
transform 1 0 25024 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _192_
timestamp 1623529830
transform -1 0 27416 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1623529830
transform 1 0 26956 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1623529830
transform -1 0 28244 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _190_
timestamp 1623529830
transform 1 0 28244 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _242_
timestamp 1623529830
transform 1 0 28612 0 1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1623529830
transform 1 0 27784 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1623529830
transform 1 0 27324 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1623529830
transform 1 0 27416 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_291
timestamp 1623529830
transform 1 0 27876 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_286
timestamp 1623529830
transform 1 0 27416 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_295
timestamp 1623529830
transform 1 0 28244 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _176_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform -1 0 31648 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _194_
timestamp 1623529830
transform -1 0 32752 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1623529830
transform 1 0 30452 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_315
timestamp 1623529830
transform 1 0 30084 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_320
timestamp 1623529830
transform 1 0 30544 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_320
timestamp 1623529830
transform 1 0 30544 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _232_
timestamp 1623529830
transform -1 0 34868 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1623529830
transform 1 0 33120 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1623529830
transform 1 0 32568 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_344
timestamp 1623529830
transform 1 0 32752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1623529830
transform 1 0 33212 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_332
timestamp 1623529830
transform 1 0 31648 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_340
timestamp 1623529830
transform 1 0 32384 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_343
timestamp 1623529830
transform 1 0 32660 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _177_
timestamp 1623529830
transform 1 0 35236 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _243_
timestamp 1623529830
transform 1 0 33580 0 -1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_1_367
timestamp 1623529830
transform 1 0 34868 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_379
timestamp 1623529830
transform 1 0 35972 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_378
timestamp 1623529830
transform 1 0 35880 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_373
timestamp 1623529830
transform 1 0 35420 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1623529830
transform 1 0 35788 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_386
timestamp 1623529830
transform 1 0 36616 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output4
timestamp 1623529830
transform -1 0 36616 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _175_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform -1 0 36984 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_1_390
timestamp 1623529830
transform 1 0 36984 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_393
timestamp 1623529830
transform 1 0 37260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _142_
timestamp 1623529830
transform 1 0 36984 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _150_
timestamp 1623529830
transform 1 0 37628 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1623529830
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1623529830
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1623529830
transform 1 0 38456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1623529830
transform 1 0 37812 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_400
timestamp 1623529830
transform 1 0 37904 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_398
timestamp 1623529830
transform 1 0 37720 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_400
timestamp 1623529830
transform 1 0 37904 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_406
timestamp 1623529830
transform 1 0 38456 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1623529830
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1623529830
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1623529830
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1623529830
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1623529830
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_30
timestamp 1623529830
transform 1 0 3864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_42
timestamp 1623529830
transform 1 0 4968 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_54
timestamp 1623529830
transform 1 0 6072 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1623529830
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_66
timestamp 1623529830
transform 1 0 7176 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_78
timestamp 1623529830
transform 1 0 8280 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_87
timestamp 1623529830
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_99
timestamp 1623529830
transform 1 0 10212 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_111
timestamp 1623529830
transform 1 0 11316 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1623529830
transform 1 0 12420 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _233_
timestamp 1623529830
transform 1 0 15088 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1623529830
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_135
timestamp 1623529830
transform 1 0 13524 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_144
timestamp 1623529830
transform 1 0 14352 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_172
timestamp 1623529830
transform 1 0 16928 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _223_
timestamp 1623529830
transform 1 0 17296 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_2_196
timestamp 1623529830
transform 1 0 19136 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _206_
timestamp 1623529830
transform 1 0 20332 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1623529830
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_201
timestamp 1623529830
transform 1 0 19596 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _197_
timestamp 1623529830
transform 1 0 22540 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_2_229
timestamp 1623529830
transform 1 0 22172 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _171_
timestamp 1623529830
transform 1 0 25208 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1623529830
transform 1 0 24748 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_253
timestamp 1623529830
transform 1 0 24380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_258
timestamp 1623529830
transform 1 0 24840 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _184_
timestamp 1623529830
transform 1 0 26864 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_2_270
timestamp 1623529830
transform 1 0 25944 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_278
timestamp 1623529830
transform 1 0 26680 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _092_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform -1 0 29348 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_300
timestamp 1623529830
transform 1 0 28704 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _193_
timestamp 1623529830
transform -1 0 32292 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1623529830
transform 1 0 29992 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_307
timestamp 1623529830
transform 1 0 29348 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_313
timestamp 1623529830
transform 1 0 29900 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_315
timestamp 1623529830
transform 1 0 30084 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _227_
timestamp 1623529830
transform -1 0 34500 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_2_339
timestamp 1623529830
transform 1 0 32292 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1623529830
transform 1 0 35236 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_363
timestamp 1623529830
transform 1 0 34500 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _245_
timestamp 1623529830
transform 1 0 35696 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_2_372
timestamp 1623529830
transform 1 0 35328 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1623529830
transform 1 0 37904 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1623529830
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_396
timestamp 1623529830
transform 1 0 37536 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_403
timestamp 1623529830
transform 1 0 38180 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1623529830
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1623529830
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1623529830
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1623529830
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1623529830
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1623529830
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_51
timestamp 1623529830
transform 1 0 5796 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_58
timestamp 1623529830
transform 1 0 6440 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_70
timestamp 1623529830
transform 1 0 7544 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_82
timestamp 1623529830
transform 1 0 8648 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_94
timestamp 1623529830
transform 1 0 9752 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_106
timestamp 1623529830
transform 1 0 10856 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1623529830
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_115
timestamp 1623529830
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_127
timestamp 1623529830
transform 1 0 12788 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_139
timestamp 1623529830
transform 1 0 13892 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_151
timestamp 1623529830
transform 1 0 14996 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1623529830
transform -1 0 16468 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1623529830
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_Clk
timestamp 1623529830
transform -1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_160
timestamp 1623529830
transform 1 0 15824 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_167
timestamp 1623529830
transform 1 0 16468 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_172
timestamp 1623529830
transform 1 0 16928 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _219_
timestamp 1623529830
transform 1 0 17664 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _209_
timestamp 1623529830
transform 1 0 19872 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_3_200
timestamp 1623529830
transform 1 0 19504 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _191_
timestamp 1623529830
transform 1 0 22908 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1623529830
transform 1 0 22080 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_224
timestamp 1623529830
transform 1 0 21712 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_229
timestamp 1623529830
transform 1 0 22172 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _187_
timestamp 1623529830
transform -1 0 26956 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_3_257
timestamp 1623529830
transform 1 0 24748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_281
timestamp 1623529830
transform 1 0 26956 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _182_
timestamp 1623529830
transform 1 0 27784 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1623529830
transform 1 0 27324 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_286
timestamp 1623529830
transform 1 0 27416 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _188_
timestamp 1623529830
transform -1 0 31832 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_3_310
timestamp 1623529830
transform 1 0 29624 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _229_
timestamp 1623529830
transform -1 0 34868 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1623529830
transform 1 0 32568 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_334
timestamp 1623529830
transform 1 0 31832 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_343
timestamp 1623529830
transform 1 0 32660 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1623529830
transform 1 0 35236 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_367
timestamp 1623529830
transform 1 0 34868 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _122_
timestamp 1623529830
transform -1 0 36156 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1623529830
transform 1 0 36524 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _152_
timestamp 1623529830
transform 1 0 37168 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_374
timestamp 1623529830
transform 1 0 35512 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_381
timestamp 1623529830
transform 1 0 36156 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1623529830
transform 1 0 36800 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1623529830
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1623529830
transform 1 0 37812 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_395
timestamp 1623529830
transform 1 0 37444 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_400
timestamp 1623529830
transform 1 0 37904 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_406
timestamp 1623529830
transform 1 0 38456 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1623529830
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1623529830
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1623529830
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1623529830
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1623529830
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_30
timestamp 1623529830
transform 1 0 3864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_42
timestamp 1623529830
transform 1 0 4968 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_54
timestamp 1623529830
transform 1 0 6072 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1623529830
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_66
timestamp 1623529830
transform 1 0 7176 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_78
timestamp 1623529830
transform 1 0 8280 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_87
timestamp 1623529830
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_99
timestamp 1623529830
transform 1 0 10212 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_111
timestamp 1623529830
transform 1 0 11316 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1623529830
transform 1 0 12420 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1623529830
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_135
timestamp 1623529830
transform 1 0 13524 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_144
timestamp 1623529830
transform 1 0 14352 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1623529830
transform -1 0 16928 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_156
timestamp 1623529830
transform 1 0 15456 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_168
timestamp 1623529830
transform 1 0 16560 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_172
timestamp 1623529830
transform 1 0 16928 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _228_
timestamp 1623529830
transform 1 0 17296 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_4_196
timestamp 1623529830
transform 1 0 19136 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _212_
timestamp 1623529830
transform 1 0 20332 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1623529830
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_201
timestamp 1623529830
transform 1 0 19596 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _201_
timestamp 1623529830
transform 1 0 22540 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_4_229
timestamp 1623529830
transform 1 0 22172 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _185_
timestamp 1623529830
transform 1 0 25208 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1623529830
transform 1 0 24748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_253
timestamp 1623529830
transform 1 0 24380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_258
timestamp 1623529830
transform 1 0 24840 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_282
timestamp 1623529830
transform 1 0 27048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _180_
timestamp 1623529830
transform 1 0 27416 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _195_
timestamp 1623529830
transform 1 0 30452 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1623529830
transform 1 0 29992 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_306
timestamp 1623529830
transform 1 0 29256 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_315
timestamp 1623529830
transform 1 0 30084 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _231_
timestamp 1623529830
transform -1 0 34500 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_4_339
timestamp 1623529830
transform 1 0 32292 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1623529830
transform 1 0 35236 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_363
timestamp 1623529830
transform 1 0 34500 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1623529830
transform 1 0 35696 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 1623529830
transform 1 0 36340 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _163_
timestamp 1623529830
transform 1 0 36984 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_372
timestamp 1623529830
transform 1 0 35328 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_379
timestamp 1623529830
transform 1 0 35972 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_386
timestamp 1623529830
transform 1 0 36616 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_393
timestamp 1623529830
transform 1 0 37260 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1623529830
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_Clk
timestamp 1623529830
transform 1 0 37628 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_400
timestamp 1623529830
transform 1 0 37904 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_406
timestamp 1623529830
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1623529830
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1623529830
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1623529830
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1623529830
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1623529830
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1623529830
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_51
timestamp 1623529830
transform 1 0 5796 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_58
timestamp 1623529830
transform 1 0 6440 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_70
timestamp 1623529830
transform 1 0 7544 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_82
timestamp 1623529830
transform 1 0 8648 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_94
timestamp 1623529830
transform 1 0 9752 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_106
timestamp 1623529830
transform 1 0 10856 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1623529830
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_115
timestamp 1623529830
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_127
timestamp 1623529830
transform 1 0 12788 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_139
timestamp 1623529830
transform 1 0 13892 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_151
timestamp 1623529830
transform 1 0 14996 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1623529830
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_163
timestamp 1623529830
transform 1 0 16100 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_172
timestamp 1623529830
transform 1 0 16928 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _236_
timestamp 1623529830
transform -1 0 19504 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _217_
timestamp 1623529830
transform 1 0 19872 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_5_200
timestamp 1623529830
transform 1 0 19504 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _203_
timestamp 1623529830
transform -1 0 24748 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1623529830
transform 1 0 22080 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_224
timestamp 1623529830
transform 1 0 21712 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_229
timestamp 1623529830
transform 1 0 22172 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _186_
timestamp 1623529830
transform 1 0 25116 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_5_257
timestamp 1623529830
transform 1 0 24748 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_281
timestamp 1623529830
transform 1 0 26956 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _181_
timestamp 1623529830
transform -1 0 29624 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1623529830
transform 1 0 27324 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_286
timestamp 1623529830
transform 1 0 27416 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _213_
timestamp 1623529830
transform 1 0 29992 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_5_310
timestamp 1623529830
transform 1 0 29624 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _246_
timestamp 1623529830
transform 1 0 33028 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1623529830
transform 1 0 32568 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_334
timestamp 1623529830
transform 1 0 31832 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_343
timestamp 1623529830
transform 1 0 32660 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1623529830
transform 1 0 35236 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_367
timestamp 1623529830
transform 1 0 34868 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1623529830
transform 1 0 35880 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1623529830
transform 1 0 36524 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_374
timestamp 1623529830
transform 1 0 35512 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_381
timestamp 1623529830
transform 1 0 36156 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_388
timestamp 1623529830
transform 1 0 36800 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1623529830
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1623529830
transform 1 0 37812 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_396
timestamp 1623529830
transform 1 0 37536 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_400
timestamp 1623529830
transform 1 0 37904 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_406
timestamp 1623529830
transform 1 0 38456 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1623529830
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1623529830
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1623529830
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1623529830
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1623529830
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1623529830
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1623529830
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1623529830
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_30
timestamp 1623529830
transform 1 0 3864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_42
timestamp 1623529830
transform 1 0 4968 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1623529830
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1623529830
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1623529830
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_54
timestamp 1623529830
transform 1 0 6072 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_51
timestamp 1623529830
transform 1 0 5796 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_58
timestamp 1623529830
transform 1 0 6440 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1623529830
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_66
timestamp 1623529830
transform 1 0 7176 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_78
timestamp 1623529830
transform 1 0 8280 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_87
timestamp 1623529830
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_70
timestamp 1623529830
transform 1 0 7544 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_82
timestamp 1623529830
transform 1 0 8648 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_99
timestamp 1623529830
transform 1 0 10212 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_94
timestamp 1623529830
transform 1 0 9752 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_106
timestamp 1623529830
transform 1 0 10856 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1623529830
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_111
timestamp 1623529830
transform 1 0 11316 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_123
timestamp 1623529830
transform 1 0 12420 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_115
timestamp 1623529830
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_127
timestamp 1623529830
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1623529830
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_135
timestamp 1623529830
transform 1 0 13524 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_144
timestamp 1623529830
transform 1 0 14352 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_139
timestamp 1623529830
transform 1 0 13892 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_151
timestamp 1623529830
transform 1 0 14996 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1623529830
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_156
timestamp 1623529830
transform 1 0 15456 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_168
timestamp 1623529830
transform 1 0 16560 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_163
timestamp 1623529830
transform 1 0 16100 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_172
timestamp 1623529830
transform 1 0 16928 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _110_
timestamp 1623529830
transform -1 0 19136 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1623529830
transform -1 0 18492 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_Clk
timestamp 1623529830
transform 1 0 17388 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_176
timestamp 1623529830
transform 1 0 17296 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_180
timestamp 1623529830
transform 1 0 17664 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_189
timestamp 1623529830
transform 1 0 18492 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_196
timestamp 1623529830
transform 1 0 19136 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1623529830
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_196
timestamp 1623529830
transform 1 0 19136 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1623529830
transform 1 0 19228 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _218_
timestamp 1623529830
transform 1 0 20332 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _222_
timestamp 1623529830
transform 1 0 19872 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1623529830
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_201
timestamp 1623529830
transform 1 0 19596 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_200
timestamp 1623529830
transform 1 0 19504 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _208_
timestamp 1623529830
transform 1 0 22540 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _211_
timestamp 1623529830
transform 1 0 22908 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1623529830
transform 1 0 22080 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_229
timestamp 1623529830
transform 1 0 22172 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_224
timestamp 1623529830
transform 1 0 21712 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_229
timestamp 1623529830
transform 1 0 22172 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _172_
timestamp 1623529830
transform 1 0 25208 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _199_
timestamp 1623529830
transform 1 0 25116 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1623529830
transform 1 0 24748 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_253
timestamp 1623529830
transform 1 0 24380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_258
timestamp 1623529830
transform 1 0 24840 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_257
timestamp 1623529830
transform 1 0 24748 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _097_
timestamp 1623529830
transform -1 0 26588 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _183_
timestamp 1623529830
transform -1 0 28796 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_6_270
timestamp 1623529830
transform 1 0 25944 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_277
timestamp 1623529830
transform 1 0 26588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_281
timestamp 1623529830
transform 1 0 26956 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _091_
timestamp 1623529830
transform 1 0 29164 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _196_
timestamp 1623529830
transform 1 0 27784 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1623529830
transform 1 0 27324 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_301
timestamp 1623529830
transform 1 0 28796 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_286
timestamp 1623529830
transform 1 0 27416 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _221_
timestamp 1623529830
transform -1 0 32292 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _230_
timestamp 1623529830
transform -1 0 31832 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1623529830
transform 1 0 29992 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_308
timestamp 1623529830
transform 1 0 29440 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_315
timestamp 1623529830
transform 1 0 30084 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_310
timestamp 1623529830
transform 1 0 29624 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1623529830
transform 1 0 32660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1623529830
transform 1 0 33028 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1623529830
transform 1 0 32568 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_339
timestamp 1623529830
transform 1 0 32292 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_346
timestamp 1623529830
transform 1 0 32936 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_334
timestamp 1623529830
transform 1 0 31832 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_343
timestamp 1623529830
transform 1 0 32660 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_357
timestamp 1623529830
transform 1 0 33948 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_350
timestamp 1623529830
transform 1 0 33304 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_360
timestamp 1623529830
transform 1 0 34224 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_353
timestamp 1623529830
transform 1 0 33580 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 1623529830
transform 1 0 33672 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _128_
timestamp 1623529830
transform -1 0 34224 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1623529830
transform 1 0 33304 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_364
timestamp 1623529830
transform 1 0 34592 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_367
timestamp 1623529830
transform 1 0 34868 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1623529830
transform 1 0 35236 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1623529830
transform 1 0 34960 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _157_
timestamp 1623529830
transform 1 0 34316 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp 1623529830
transform 1 0 34592 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_371
timestamp 1623529830
transform 1 0 35236 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1623529830
transform 1 0 35696 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_372
timestamp 1623529830
transform 1 0 35328 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_379
timestamp 1623529830
transform 1 0 35972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_391
timestamp 1623529830
transform 1 0 37076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_383
timestamp 1623529830
transform 1 0 36340 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1623529830
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1623529830
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1623529830
transform 1 0 37812 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_403
timestamp 1623529830
transform 1 0 38180 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_395
timestamp 1623529830
transform 1 0 37444 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_400
timestamp 1623529830
transform 1 0 37904 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_406
timestamp 1623529830
transform 1 0 38456 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1623529830
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1623529830
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1623529830
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1623529830
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1623529830
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_30
timestamp 1623529830
transform 1 0 3864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_42
timestamp 1623529830
transform 1 0 4968 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_54
timestamp 1623529830
transform 1 0 6072 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1623529830
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_66
timestamp 1623529830
transform 1 0 7176 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_78
timestamp 1623529830
transform 1 0 8280 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_87
timestamp 1623529830
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_99
timestamp 1623529830
transform 1 0 10212 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_111
timestamp 1623529830
transform 1 0 11316 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1623529830
transform 1 0 12420 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1623529830
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_135
timestamp 1623529830
transform 1 0 13524 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_144
timestamp 1623529830
transform 1 0 14352 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_156
timestamp 1623529830
transform 1 0 15456 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_168
timestamp 1623529830
transform 1 0 16560 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_180
timestamp 1623529830
transform 1 0 17664 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_192
timestamp 1623529830
transform 1 0 18768 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _234_
timestamp 1623529830
transform 1 0 20332 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1623529830
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_201
timestamp 1623529830
transform 1 0 19596 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _215_
timestamp 1623529830
transform 1 0 22540 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_8_229
timestamp 1623529830
transform 1 0 22172 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1623529830
transform 1 0 24748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_253
timestamp 1623529830
transform 1 0 24380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_258
timestamp 1623529830
transform 1 0 24840 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _098_
timestamp 1623529830
transform 1 0 25668 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _198_
timestamp 1623529830
transform -1 0 28152 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_8_266
timestamp 1623529830
transform 1 0 25576 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_270
timestamp 1623529830
transform 1 0 25944 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1623529830
transform -1 0 28888 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_294
timestamp 1623529830
transform 1 0 28152 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_298
timestamp 1623529830
transform 1 0 28520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_302
timestamp 1623529830
transform 1 0 28888 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1623529830
transform -1 0 29532 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _244_
timestamp 1623529830
transform -1 0 32292 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1623529830
transform 1 0 29992 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_309
timestamp 1623529830
transform 1 0 29532 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_313
timestamp 1623529830
transform 1 0 29900 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_315
timestamp 1623529830
transform 1 0 30084 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _147_
timestamp 1623529830
transform 1 0 32660 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_339
timestamp 1623529830
transform 1 0 32292 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_346
timestamp 1623529830
transform 1 0 32936 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _153_
timestamp 1623529830
transform 1 0 33304 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1623529830
transform 1 0 33948 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1623529830
transform 1 0 35236 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_Clk
timestamp 1623529830
transform -1 0 34868 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_353
timestamp 1623529830
transform 1 0 33580 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_360
timestamp 1623529830
transform 1 0 34224 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_367
timestamp 1623529830
transform 1 0 34868 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_372
timestamp 1623529830
transform 1 0 35328 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_384
timestamp 1623529830
transform 1 0 36432 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1623529830
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_396
timestamp 1623529830
transform 1 0 37536 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_404
timestamp 1623529830
transform 1 0 38272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1623529830
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1623529830
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1623529830
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1623529830
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1623529830
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1623529830
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_51
timestamp 1623529830
transform 1 0 5796 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_58
timestamp 1623529830
transform 1 0 6440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_70
timestamp 1623529830
transform 1 0 7544 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_82
timestamp 1623529830
transform 1 0 8648 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_94
timestamp 1623529830
transform 1 0 9752 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_106
timestamp 1623529830
transform 1 0 10856 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1623529830
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_115
timestamp 1623529830
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_127
timestamp 1623529830
transform 1 0 12788 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_139
timestamp 1623529830
transform 1 0 13892 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_151
timestamp 1623529830
transform 1 0 14996 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1623529830
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_163
timestamp 1623529830
transform 1 0 16100 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_172
timestamp 1623529830
transform 1 0 16928 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1623529830
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_196
timestamp 1623529830
transform 1 0 19136 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1623529830
transform 1 0 20792 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_Clk
timestamp 1623529830
transform 1 0 20056 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_204
timestamp 1623529830
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_209
timestamp 1623529830
transform 1 0 20332 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_213
timestamp 1623529830
transform 1 0 20700 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_217
timestamp 1623529830
transform 1 0 21068 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1623529830
transform -1 0 21712 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _170_
timestamp 1623529830
transform 1 0 23092 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1623529830
transform 1 0 22080 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_224
timestamp 1623529830
transform 1 0 21712 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_229
timestamp 1623529830
transform 1 0 22172 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_237
timestamp 1623529830
transform 1 0 22908 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _207_
timestamp 1623529830
transform 1 0 24564 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_9_246
timestamp 1623529830
transform 1 0 23736 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_254
timestamp 1623529830
transform 1 0 24472 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_275
timestamp 1623529830
transform 1 0 26404 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_283
timestamp 1623529830
transform 1 0 27140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_1  _216_
timestamp 1623529830
transform -1 0 29624 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1623529830
transform 1 0 27324 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_286
timestamp 1623529830
transform 1 0 27416 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1623529830
transform -1 0 30268 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1623529830
transform 1 0 30636 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_310
timestamp 1623529830
transform 1 0 29624 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_317
timestamp 1623529830
transform 1 0 30268 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_324
timestamp 1623529830
transform 1 0 30912 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1623529830
transform 1 0 31280 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _143_
timestamp 1623529830
transform 1 0 31924 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1623529830
transform 1 0 33028 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1623529830
transform 1 0 32568 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_331
timestamp 1623529830
transform 1 0 31556 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_338
timestamp 1623529830
transform 1 0 32200 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_343
timestamp 1623529830
transform 1 0 32660 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1623529830
transform -1 0 33948 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_350
timestamp 1623529830
transform 1 0 33304 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_357
timestamp 1623529830
transform 1 0 33948 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_369
timestamp 1623529830
transform 1 0 35052 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_381
timestamp 1623529830
transform 1 0 36156 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_393
timestamp 1623529830
transform 1 0 37260 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1623529830
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1623529830
transform 1 0 37812 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_400
timestamp 1623529830
transform 1 0 37904 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_406
timestamp 1623529830
transform 1 0 38456 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1623529830
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1623529830
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1623529830
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1623529830
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1623529830
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1623529830
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1623529830
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_54
timestamp 1623529830
transform 1 0 6072 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1623529830
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_66
timestamp 1623529830
transform 1 0 7176 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_78
timestamp 1623529830
transform 1 0 8280 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_87
timestamp 1623529830
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_99
timestamp 1623529830
transform 1 0 10212 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_111
timestamp 1623529830
transform 1 0 11316 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1623529830
transform 1 0 12420 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1623529830
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_135
timestamp 1623529830
transform 1 0 13524 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_144
timestamp 1623529830
transform 1 0 14352 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_156
timestamp 1623529830
transform 1 0 15456 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_168
timestamp 1623529830
transform 1 0 16560 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_180
timestamp 1623529830
transform 1 0 17664 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_192
timestamp 1623529830
transform 1 0 18768 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1623529830
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_201
timestamp 1623529830
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_213
timestamp 1623529830
transform 1 0 20700 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1623529830
transform 1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _225_
timestamp 1623529830
transform -1 0 24380 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_Clk
timestamp 1623529830
transform -1 0 21528 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_222
timestamp 1623529830
transform 1 0 21528 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_229
timestamp 1623529830
transform 1 0 22172 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _210_
timestamp 1623529830
transform 1 0 25208 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1623529830
transform 1 0 24748 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_253
timestamp 1623529830
transform 1 0 24380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_258
timestamp 1623529830
transform 1 0 24840 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_282
timestamp 1623529830
transform 1 0 27048 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _247_
timestamp 1623529830
transform 1 0 27784 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1623529830
transform 1 0 30452 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _144_
timestamp 1623529830
transform 1 0 31096 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1623529830
transform 1 0 29992 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_310
timestamp 1623529830
transform 1 0 29624 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_315
timestamp 1623529830
transform 1 0 30084 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_322
timestamp 1623529830
transform 1 0 30728 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _156_
timestamp 1623529830
transform 1 0 31740 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1623529830
transform 1 0 32384 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_Clk
timestamp 1623529830
transform 1 0 33028 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_329
timestamp 1623529830
transform 1 0 31372 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_336
timestamp 1623529830
transform 1 0 32016 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_343
timestamp 1623529830
transform 1 0 32660 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1623529830
transform 1 0 35236 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_350
timestamp 1623529830
transform 1 0 33304 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_362
timestamp 1623529830
transform 1 0 34408 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_370
timestamp 1623529830
transform 1 0 35144 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_372
timestamp 1623529830
transform 1 0 35328 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_384
timestamp 1623529830
transform 1 0 36432 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1623529830
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_396
timestamp 1623529830
transform 1 0 37536 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_404
timestamp 1623529830
transform 1 0 38272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1623529830
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1623529830
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1623529830
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1623529830
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1623529830
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1623529830
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_51
timestamp 1623529830
transform 1 0 5796 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_58
timestamp 1623529830
transform 1 0 6440 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_70
timestamp 1623529830
transform 1 0 7544 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_82
timestamp 1623529830
transform 1 0 8648 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_94
timestamp 1623529830
transform 1 0 9752 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_106
timestamp 1623529830
transform 1 0 10856 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1623529830
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_115
timestamp 1623529830
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_127
timestamp 1623529830
transform 1 0 12788 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_139
timestamp 1623529830
transform 1 0 13892 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_151
timestamp 1623529830
transform 1 0 14996 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1623529830
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_163
timestamp 1623529830
transform 1 0 16100 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_172
timestamp 1623529830
transform 1 0 16928 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1623529830
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1623529830
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1623529830
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1623529830
transform -1 0 23092 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1623529830
transform 1 0 22080 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_220
timestamp 1623529830
transform 1 0 21344 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_229
timestamp 1623529830
transform 1 0 22172 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_235
timestamp 1623529830
transform 1 0 22724 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_239
timestamp 1623529830
transform 1 0 23092 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1623529830
transform 1 0 24104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1623529830
transform 1 0 23460 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _214_
timestamp 1623529830
transform 1 0 25116 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_11_246
timestamp 1623529830
transform 1 0 23736 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_253
timestamp 1623529830
transform 1 0 24380 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_281
timestamp 1623529830
transform 1 0 26956 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _248_
timestamp 1623529830
transform -1 0 29624 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1623529830
transform 1 0 27324 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_286
timestamp 1623529830
transform 1 0 27416 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _090_
timestamp 1623529830
transform -1 0 31464 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _129_
timestamp 1623529830
transform 1 0 29992 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_310
timestamp 1623529830
transform 1 0 29624 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_317
timestamp 1623529830
transform 1 0 30268 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_325
timestamp 1623529830
transform 1 0 31004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1623529830
transform 1 0 31832 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1623529830
transform 1 0 32568 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_330
timestamp 1623529830
transform 1 0 31464 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_337
timestamp 1623529830
transform 1 0 32108 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_341
timestamp 1623529830
transform 1 0 32476 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_343
timestamp 1623529830
transform 1 0 32660 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_355
timestamp 1623529830
transform 1 0 33764 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_367
timestamp 1623529830
transform 1 0 34868 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_379
timestamp 1623529830
transform 1 0 35972 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_391
timestamp 1623529830
transform 1 0 37076 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1623529830
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1623529830
transform 1 0 37812 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_400
timestamp 1623529830
transform 1 0 37904 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_406
timestamp 1623529830
transform 1 0 38456 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1623529830
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1623529830
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1623529830
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1623529830
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1623529830
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_30
timestamp 1623529830
transform 1 0 3864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_42
timestamp 1623529830
transform 1 0 4968 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_54
timestamp 1623529830
transform 1 0 6072 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1623529830
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_66
timestamp 1623529830
transform 1 0 7176 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_78
timestamp 1623529830
transform 1 0 8280 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_87
timestamp 1623529830
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_99
timestamp 1623529830
transform 1 0 10212 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_111
timestamp 1623529830
transform 1 0 11316 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_123
timestamp 1623529830
transform 1 0 12420 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1623529830
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_135
timestamp 1623529830
transform 1 0 13524 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_144
timestamp 1623529830
transform 1 0 14352 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_156
timestamp 1623529830
transform 1 0 15456 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_168
timestamp 1623529830
transform 1 0 16560 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_180
timestamp 1623529830
transform 1 0 17664 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_192
timestamp 1623529830
transform 1 0 18768 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1623529830
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_201
timestamp 1623529830
transform 1 0 19596 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_213
timestamp 1623529830
transform 1 0 20700 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_Clk
timestamp 1623529830
transform 1 0 22816 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_225
timestamp 1623529830
transform 1 0 21804 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_233
timestamp 1623529830
transform 1 0 22540 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_239
timestamp 1623529830
transform 1 0 23092 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1623529830
transform -1 0 24380 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 1623529830
transform 1 0 23460 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _220_
timestamp 1623529830
transform -1 0 27048 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1623529830
transform 1 0 24748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_246
timestamp 1623529830
transform 1 0 23736 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_253
timestamp 1623529830
transform 1 0 24380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_258
timestamp 1623529830
transform 1 0 24840 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_282
timestamp 1623529830
transform 1 0 27048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _116_
timestamp 1623529830
transform 1 0 27416 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1623529830
transform -1 0 28336 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1623529830
transform 1 0 28704 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_289
timestamp 1623529830
transform 1 0 27692 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_296
timestamp 1623529830
transform 1 0 28336 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_303
timestamp 1623529830
transform 1 0 28980 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 1623529830
transform 1 0 29348 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1623529830
transform 1 0 30452 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1623529830
transform 1 0 29992 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_Clk
timestamp 1623529830
transform 1 0 31096 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_310
timestamp 1623529830
transform 1 0 29624 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_315
timestamp 1623529830
transform 1 0 30084 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_322
timestamp 1623529830
transform 1 0 30728 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_329
timestamp 1623529830
transform 1 0 31372 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_341
timestamp 1623529830
transform 1 0 32476 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1623529830
transform 1 0 35236 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_353
timestamp 1623529830
transform 1 0 33580 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_365
timestamp 1623529830
transform 1 0 34684 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_372
timestamp 1623529830
transform 1 0 35328 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_384
timestamp 1623529830
transform 1 0 36432 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1623529830
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_396
timestamp 1623529830
transform 1 0 37536 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_404
timestamp 1623529830
transform 1 0 38272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1623529830
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1623529830
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1623529830
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1623529830
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1623529830
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1623529830
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1623529830
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1623529830
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1623529830
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1623529830
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1623529830
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_42
timestamp 1623529830
transform 1 0 4968 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1623529830
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_51
timestamp 1623529830
transform 1 0 5796 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_58
timestamp 1623529830
transform 1 0 6440 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_54
timestamp 1623529830
transform 1 0 6072 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1623529830
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_70
timestamp 1623529830
transform 1 0 7544 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_82
timestamp 1623529830
transform 1 0 8648 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_66
timestamp 1623529830
transform 1 0 7176 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_78
timestamp 1623529830
transform 1 0 8280 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_87
timestamp 1623529830
transform 1 0 9108 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_94
timestamp 1623529830
transform 1 0 9752 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_106
timestamp 1623529830
transform 1 0 10856 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_99
timestamp 1623529830
transform 1 0 10212 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1623529830
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_115
timestamp 1623529830
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_127
timestamp 1623529830
transform 1 0 12788 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_111
timestamp 1623529830
transform 1 0 11316 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_123
timestamp 1623529830
transform 1 0 12420 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1623529830
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_139
timestamp 1623529830
transform 1 0 13892 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_151
timestamp 1623529830
transform 1 0 14996 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_135
timestamp 1623529830
transform 1 0 13524 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_144
timestamp 1623529830
transform 1 0 14352 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1623529830
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_163
timestamp 1623529830
transform 1 0 16100 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_172
timestamp 1623529830
transform 1 0 16928 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_156
timestamp 1623529830
transform 1 0 15456 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_168
timestamp 1623529830
transform 1 0 16560 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1623529830
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1623529830
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_180
timestamp 1623529830
transform 1 0 17664 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_192
timestamp 1623529830
transform 1 0 18768 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1623529830
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1623529830
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_201
timestamp 1623529830
transform 1 0 19596 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_213
timestamp 1623529830
transform 1 0 20700 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1623529830
transform 1 0 22080 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_220
timestamp 1623529830
transform 1 0 21344 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_229
timestamp 1623529830
transform 1 0 22172 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_225
timestamp 1623529830
transform 1 0 21804 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_237
timestamp 1623529830
transform 1 0 22908 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_249
timestamp 1623529830
transform 1 0 24012 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_250
timestamp 1623529830
transform 1 0 24104 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_241
timestamp 1623529830
transform 1 0 23276 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_Clk
timestamp 1623529830
transform -1 0 24380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1623529830
transform 1 0 23828 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_258
timestamp 1623529830
transform 1 0 24840 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_253
timestamp 1623529830
transform 1 0 24380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_257
timestamp 1623529830
transform 1 0 24748 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1623529830
transform 1 0 24748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1623529830
transform 1 0 24472 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_Clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform 1 0 25116 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1623529830
transform 1 0 25760 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1623529830
transform 1 0 26404 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1623529830
transform 1 0 27048 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_281
timestamp 1623529830
transform 1 0 26956 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_266
timestamp 1623529830
transform 1 0 25576 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_271
timestamp 1623529830
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_278
timestamp 1623529830
transform 1 0 26680 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_285
timestamp 1623529830
transform 1 0 27324 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_286
timestamp 1623529830
transform 1 0 27416 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1623529830
transform 1 0 27324 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_292
timestamp 1623529830
transform 1 0 27968 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_293
timestamp 1623529830
transform 1 0 28060 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _141_
timestamp 1623529830
transform 1 0 27692 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _104_
timestamp 1623529830
transform -1 0 28060 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1623529830
transform 1 0 28336 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1623529830
transform 1 0 28428 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_299
timestamp 1623529830
transform 1 0 28612 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_300
timestamp 1623529830
transform 1 0 28704 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _159_
timestamp 1623529830
transform 1 0 28980 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _145_
timestamp 1623529830
transform 1 0 29072 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_315
timestamp 1623529830
transform 1 0 30084 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_306
timestamp 1623529830
transform 1 0 29256 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_314
timestamp 1623529830
transform 1 0 29992 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_307
timestamp 1623529830
transform 1 0 29348 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1623529830
transform 1 0 29992 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1623529830
transform 1 0 29716 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_Clk
timestamp 1623529830
transform -1 0 31096 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1623529830
transform 1 0 30360 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_326
timestamp 1623529830
transform 1 0 31096 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_321
timestamp 1623529830
transform 1 0 30636 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1623529830
transform 1 0 32568 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_333
timestamp 1623529830
transform 1 0 31740 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_341
timestamp 1623529830
transform 1 0 32476 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_343
timestamp 1623529830
transform 1 0 32660 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_338
timestamp 1623529830
transform 1 0 32200 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1623529830
transform 1 0 35236 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_355
timestamp 1623529830
transform 1 0 33764 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_367
timestamp 1623529830
transform 1 0 34868 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_350
timestamp 1623529830
transform 1 0 33304 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_362
timestamp 1623529830
transform 1 0 34408 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_370
timestamp 1623529830
transform 1 0 35144 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_379
timestamp 1623529830
transform 1 0 35972 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_391
timestamp 1623529830
transform 1 0 37076 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_372
timestamp 1623529830
transform 1 0 35328 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_384
timestamp 1623529830
transform 1 0 36432 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1623529830
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1623529830
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1623529830
transform 1 0 37812 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_400
timestamp 1623529830
transform 1 0 37904 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_406
timestamp 1623529830
transform 1 0 38456 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_396
timestamp 1623529830
transform 1 0 37536 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_404
timestamp 1623529830
transform 1 0 38272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1623529830
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1623529830
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1623529830
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1623529830
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1623529830
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1623529830
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_51
timestamp 1623529830
transform 1 0 5796 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_58
timestamp 1623529830
transform 1 0 6440 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_70
timestamp 1623529830
transform 1 0 7544 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_82
timestamp 1623529830
transform 1 0 8648 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_94
timestamp 1623529830
transform 1 0 9752 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_106
timestamp 1623529830
transform 1 0 10856 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1623529830
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_115
timestamp 1623529830
transform 1 0 11684 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_127
timestamp 1623529830
transform 1 0 12788 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_139
timestamp 1623529830
transform 1 0 13892 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_151
timestamp 1623529830
transform 1 0 14996 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1623529830
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_163
timestamp 1623529830
transform 1 0 16100 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_172
timestamp 1623529830
transform 1 0 16928 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1623529830
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1623529830
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1623529830
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1623529830
transform 1 0 22080 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_220
timestamp 1623529830
transform 1 0 21344 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_229
timestamp 1623529830
transform 1 0 22172 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_241
timestamp 1623529830
transform 1 0 23276 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_253
timestamp 1623529830
transform 1 0 24380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1623529830
transform -1 0 25760 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 1623529830
transform 1 0 26128 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_268
timestamp 1623529830
transform 1 0 25760 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_275
timestamp 1623529830
transform 1 0 26404 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_283
timestamp 1623529830
transform 1 0 27140 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1623529830
transform 1 0 27324 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_Clk
timestamp 1623529830
transform 1 0 27784 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_286
timestamp 1623529830
transform 1 0 27416 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1623529830
transform 1 0 28060 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1623529830
transform 1 0 29164 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1623529830
transform 1 0 30268 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1623529830
transform 1 0 32568 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_329
timestamp 1623529830
transform 1 0 31372 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_341
timestamp 1623529830
transform 1 0 32476 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_343
timestamp 1623529830
transform 1 0 32660 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_355
timestamp 1623529830
transform 1 0 33764 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_367
timestamp 1623529830
transform 1 0 34868 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_379
timestamp 1623529830
transform 1 0 35972 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_391
timestamp 1623529830
transform 1 0 37076 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1623529830
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1623529830
transform 1 0 37812 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_400
timestamp 1623529830
transform 1 0 37904 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_406
timestamp 1623529830
transform 1 0 38456 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1623529830
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1623529830
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1623529830
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1623529830
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1623529830
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_30
timestamp 1623529830
transform 1 0 3864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_42
timestamp 1623529830
transform 1 0 4968 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_54
timestamp 1623529830
transform 1 0 6072 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1623529830
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_66
timestamp 1623529830
transform 1 0 7176 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_78
timestamp 1623529830
transform 1 0 8280 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_87
timestamp 1623529830
transform 1 0 9108 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_99
timestamp 1623529830
transform 1 0 10212 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_111
timestamp 1623529830
transform 1 0 11316 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_123
timestamp 1623529830
transform 1 0 12420 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1623529830
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_135
timestamp 1623529830
transform 1 0 13524 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_144
timestamp 1623529830
transform 1 0 14352 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_156
timestamp 1623529830
transform 1 0 15456 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_168
timestamp 1623529830
transform 1 0 16560 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_180
timestamp 1623529830
transform 1 0 17664 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_192
timestamp 1623529830
transform 1 0 18768 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1623529830
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_201
timestamp 1623529830
transform 1 0 19596 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_213
timestamp 1623529830
transform 1 0 20700 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_225
timestamp 1623529830
transform 1 0 21804 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_237
timestamp 1623529830
transform 1 0 22908 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1623529830
transform 1 0 24748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_249
timestamp 1623529830
transform 1 0 24012 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_258
timestamp 1623529830
transform 1 0 24840 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _135_
timestamp 1623529830
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_270
timestamp 1623529830
transform 1 0 25944 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1623529830
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_280
timestamp 1623529830
transform 1 0 26864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_292
timestamp 1623529830
transform 1 0 27968 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_304
timestamp 1623529830
transform 1 0 29072 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1623529830
transform 1 0 29992 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_312
timestamp 1623529830
transform 1 0 29808 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_315
timestamp 1623529830
transform 1 0 30084 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_327
timestamp 1623529830
transform 1 0 31188 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _237_
timestamp 1623529830
transform -1 0 33488 0 -1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1623529830
transform 1 0 35236 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_352
timestamp 1623529830
transform 1 0 33488 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_364
timestamp 1623529830
transform 1 0 34592 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_370
timestamp 1623529830
transform 1 0 35144 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_372
timestamp 1623529830
transform 1 0 35328 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_384
timestamp 1623529830
transform 1 0 36432 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1623529830
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_396
timestamp 1623529830
transform 1 0 37536 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_404
timestamp 1623529830
transform 1 0 38272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1623529830
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1623529830
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1623529830
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1623529830
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1623529830
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1623529830
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_51
timestamp 1623529830
transform 1 0 5796 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_58
timestamp 1623529830
transform 1 0 6440 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_70
timestamp 1623529830
transform 1 0 7544 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_82
timestamp 1623529830
transform 1 0 8648 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_94
timestamp 1623529830
transform 1 0 9752 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_106
timestamp 1623529830
transform 1 0 10856 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1623529830
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_115
timestamp 1623529830
transform 1 0 11684 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_127
timestamp 1623529830
transform 1 0 12788 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_139
timestamp 1623529830
transform 1 0 13892 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_151
timestamp 1623529830
transform 1 0 14996 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1623529830
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_163
timestamp 1623529830
transform 1 0 16100 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_172
timestamp 1623529830
transform 1 0 16928 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1623529830
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1623529830
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1623529830
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1623529830
transform 1 0 22080 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_220
timestamp 1623529830
transform 1 0 21344 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_229
timestamp 1623529830
transform 1 0 22172 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_241
timestamp 1623529830
transform 1 0 23276 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_253
timestamp 1623529830
transform 1 0 24380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_265
timestamp 1623529830
transform 1 0 25484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_277
timestamp 1623529830
transform 1 0 26588 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1623529830
transform 1 0 27324 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_286
timestamp 1623529830
transform 1 0 27416 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_298
timestamp 1623529830
transform 1 0 28520 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_310
timestamp 1623529830
transform 1 0 29624 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_322
timestamp 1623529830
transform 1 0 30728 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1623529830
transform 1 0 32568 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_334
timestamp 1623529830
transform 1 0 31832 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_343
timestamp 1623529830
transform 1 0 32660 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_355
timestamp 1623529830
transform 1 0 33764 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_367
timestamp 1623529830
transform 1 0 34868 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_379
timestamp 1623529830
transform 1 0 35972 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_391
timestamp 1623529830
transform 1 0 37076 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1623529830
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1623529830
transform 1 0 37812 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_400
timestamp 1623529830
transform 1 0 37904 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_406
timestamp 1623529830
transform 1 0 38456 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1623529830
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1623529830
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1623529830
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1623529830
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1623529830
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_30
timestamp 1623529830
transform 1 0 3864 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_42
timestamp 1623529830
transform 1 0 4968 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_54
timestamp 1623529830
transform 1 0 6072 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1623529830
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_66
timestamp 1623529830
transform 1 0 7176 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_78
timestamp 1623529830
transform 1 0 8280 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_87
timestamp 1623529830
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_99
timestamp 1623529830
transform 1 0 10212 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_111
timestamp 1623529830
transform 1 0 11316 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_123
timestamp 1623529830
transform 1 0 12420 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1623529830
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_135
timestamp 1623529830
transform 1 0 13524 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_144
timestamp 1623529830
transform 1 0 14352 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_156
timestamp 1623529830
transform 1 0 15456 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_168
timestamp 1623529830
transform 1 0 16560 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_180
timestamp 1623529830
transform 1 0 17664 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_192
timestamp 1623529830
transform 1 0 18768 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1623529830
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_201
timestamp 1623529830
transform 1 0 19596 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_213
timestamp 1623529830
transform 1 0 20700 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_225
timestamp 1623529830
transform 1 0 21804 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_237
timestamp 1623529830
transform 1 0 22908 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1623529830
transform 1 0 24748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_249
timestamp 1623529830
transform 1 0 24012 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_258
timestamp 1623529830
transform 1 0 24840 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_270
timestamp 1623529830
transform 1 0 25944 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_282
timestamp 1623529830
transform 1 0 27048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_294
timestamp 1623529830
transform 1 0 28152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _179_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform -1 0 31464 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1623529830
transform 1 0 29992 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_306
timestamp 1623529830
transform 1 0 29256 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_315
timestamp 1623529830
transform 1 0 30084 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfstp_1  _238_
timestamp 1623529830
transform 1 0 31832 0 -1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_18_330
timestamp 1623529830
transform 1 0 31464 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1623529830
transform 1 0 35236 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_355
timestamp 1623529830
transform 1 0 33764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_367
timestamp 1623529830
transform 1 0 34868 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_372
timestamp 1623529830
transform 1 0 35328 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_384
timestamp 1623529830
transform 1 0 36432 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1623529830
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_396
timestamp 1623529830
transform 1 0 37536 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_404
timestamp 1623529830
transform 1 0 38272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1623529830
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1623529830
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1623529830
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1623529830
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1623529830
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1623529830
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1623529830
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1623529830
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1623529830
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1623529830
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_30
timestamp 1623529830
transform 1 0 3864 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_42
timestamp 1623529830
transform 1 0 4968 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1623529830
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_51
timestamp 1623529830
transform 1 0 5796 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_58
timestamp 1623529830
transform 1 0 6440 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_54
timestamp 1623529830
transform 1 0 6072 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1623529830
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_70
timestamp 1623529830
transform 1 0 7544 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_82
timestamp 1623529830
transform 1 0 8648 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_66
timestamp 1623529830
transform 1 0 7176 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_78
timestamp 1623529830
transform 1 0 8280 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_87
timestamp 1623529830
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_94
timestamp 1623529830
transform 1 0 9752 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_106
timestamp 1623529830
transform 1 0 10856 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_99
timestamp 1623529830
transform 1 0 10212 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1623529830
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_115
timestamp 1623529830
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_127
timestamp 1623529830
transform 1 0 12788 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_111
timestamp 1623529830
transform 1 0 11316 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_123
timestamp 1623529830
transform 1 0 12420 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1623529830
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_139
timestamp 1623529830
transform 1 0 13892 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_151
timestamp 1623529830
transform 1 0 14996 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_135
timestamp 1623529830
transform 1 0 13524 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_144
timestamp 1623529830
transform 1 0 14352 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1623529830
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_163
timestamp 1623529830
transform 1 0 16100 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_172
timestamp 1623529830
transform 1 0 16928 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_156
timestamp 1623529830
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_168
timestamp 1623529830
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1623529830
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1623529830
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_180
timestamp 1623529830
transform 1 0 17664 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_192
timestamp 1623529830
transform 1 0 18768 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1623529830
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1623529830
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_201
timestamp 1623529830
transform 1 0 19596 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_213
timestamp 1623529830
transform 1 0 20700 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1623529830
transform 1 0 22080 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_220
timestamp 1623529830
transform 1 0 21344 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_229
timestamp 1623529830
transform 1 0 22172 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_225
timestamp 1623529830
transform 1 0 21804 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_237
timestamp 1623529830
transform 1 0 22908 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1623529830
transform 1 0 24748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_241
timestamp 1623529830
transform 1 0 23276 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_253
timestamp 1623529830
transform 1 0 24380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_249
timestamp 1623529830
transform 1 0 24012 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_258
timestamp 1623529830
transform 1 0 24840 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_265
timestamp 1623529830
transform 1 0 25484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_277
timestamp 1623529830
transform 1 0 26588 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_270
timestamp 1623529830
transform 1 0 25944 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_282
timestamp 1623529830
transform 1 0 27048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1623529830
transform 1 0 27324 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_286
timestamp 1623529830
transform 1 0 27416 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_298
timestamp 1623529830
transform 1 0 28520 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_294
timestamp 1623529830
transform 1 0 28152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfstp_1  _241_
timestamp 1623529830
transform 1 0 30268 0 1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1623529830
transform 1 0 29992 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_310
timestamp 1623529830
transform 1 0 29624 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_316
timestamp 1623529830
transform 1 0 30176 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_306
timestamp 1623529830
transform 1 0 29256 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_315
timestamp 1623529830
transform 1 0 30084 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_327
timestamp 1623529830
transform 1 0 31188 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfstp_1  _239_
timestamp 1623529830
transform -1 0 33856 0 -1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _240_
timestamp 1623529830
transform 1 0 33028 0 1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1623529830
transform 1 0 32568 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_338
timestamp 1623529830
transform 1 0 32200 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_343
timestamp 1623529830
transform 1 0 32660 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1623529830
transform 1 0 35236 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_368
timestamp 1623529830
transform 1 0 34960 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_356
timestamp 1623529830
transform 1 0 33856 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_368
timestamp 1623529830
transform 1 0 34960 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_380
timestamp 1623529830
transform 1 0 36064 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_392
timestamp 1623529830
transform 1 0 37168 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_372
timestamp 1623529830
transform 1 0 35328 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_384
timestamp 1623529830
transform 1 0 36432 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1623529830
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1623529830
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1623529830
transform 1 0 37812 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_398
timestamp 1623529830
transform 1 0 37720 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_400
timestamp 1623529830
transform 1 0 37904 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_406
timestamp 1623529830
transform 1 0 38456 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_396
timestamp 1623529830
transform 1 0 37536 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_404
timestamp 1623529830
transform 1 0 38272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1623529830
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1623529830
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1623529830
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1623529830
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1623529830
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1623529830
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_51
timestamp 1623529830
transform 1 0 5796 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_58
timestamp 1623529830
transform 1 0 6440 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_70
timestamp 1623529830
transform 1 0 7544 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_82
timestamp 1623529830
transform 1 0 8648 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_94
timestamp 1623529830
transform 1 0 9752 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_106
timestamp 1623529830
transform 1 0 10856 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1623529830
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_115
timestamp 1623529830
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_127
timestamp 1623529830
transform 1 0 12788 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_139
timestamp 1623529830
transform 1 0 13892 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_151
timestamp 1623529830
transform 1 0 14996 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1623529830
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_163
timestamp 1623529830
transform 1 0 16100 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_172
timestamp 1623529830
transform 1 0 16928 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1623529830
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1623529830
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1623529830
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1623529830
transform 1 0 22080 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_220
timestamp 1623529830
transform 1 0 21344 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_229
timestamp 1623529830
transform 1 0 22172 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_241
timestamp 1623529830
transform 1 0 23276 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_253
timestamp 1623529830
transform 1 0 24380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_265
timestamp 1623529830
transform 1 0 25484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_277
timestamp 1623529830
transform 1 0 26588 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1623529830
transform 1 0 27324 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_286
timestamp 1623529830
transform 1 0 27416 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_298
timestamp 1623529830
transform 1 0 28520 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_310
timestamp 1623529830
transform 1 0 29624 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_322
timestamp 1623529830
transform 1 0 30728 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1623529830
transform 1 0 32568 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_334
timestamp 1623529830
transform 1 0 31832 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_343
timestamp 1623529830
transform 1 0 32660 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_355
timestamp 1623529830
transform 1 0 33764 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_367
timestamp 1623529830
transform 1 0 34868 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_379
timestamp 1623529830
transform 1 0 35972 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_391
timestamp 1623529830
transform 1 0 37076 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1623529830
transform -1 0 38824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1623529830
transform 1 0 37812 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_400
timestamp 1623529830
transform 1 0 37904 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_406
timestamp 1623529830
transform 1 0 38456 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1623529830
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1623529830
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1623529830
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1623529830
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1623529830
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_30
timestamp 1623529830
transform 1 0 3864 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_42
timestamp 1623529830
transform 1 0 4968 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_54
timestamp 1623529830
transform 1 0 6072 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1623529830
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_66
timestamp 1623529830
transform 1 0 7176 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_78
timestamp 1623529830
transform 1 0 8280 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_87
timestamp 1623529830
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_99
timestamp 1623529830
transform 1 0 10212 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_111
timestamp 1623529830
transform 1 0 11316 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_123
timestamp 1623529830
transform 1 0 12420 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1623529830
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_135
timestamp 1623529830
transform 1 0 13524 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_144
timestamp 1623529830
transform 1 0 14352 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_156
timestamp 1623529830
transform 1 0 15456 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_168
timestamp 1623529830
transform 1 0 16560 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_180
timestamp 1623529830
transform 1 0 17664 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_192
timestamp 1623529830
transform 1 0 18768 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1623529830
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_201
timestamp 1623529830
transform 1 0 19596 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_213
timestamp 1623529830
transform 1 0 20700 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_225
timestamp 1623529830
transform 1 0 21804 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_237
timestamp 1623529830
transform 1 0 22908 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1623529830
transform 1 0 24748 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_249
timestamp 1623529830
transform 1 0 24012 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_258
timestamp 1623529830
transform 1 0 24840 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_270
timestamp 1623529830
transform 1 0 25944 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_282
timestamp 1623529830
transform 1 0 27048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_294
timestamp 1623529830
transform 1 0 28152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1623529830
transform 1 0 29992 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_306
timestamp 1623529830
transform 1 0 29256 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_315
timestamp 1623529830
transform 1 0 30084 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_327
timestamp 1623529830
transform 1 0 31188 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_339
timestamp 1623529830
transform 1 0 32292 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1623529830
transform 1 0 35236 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_351
timestamp 1623529830
transform 1 0 33396 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_363
timestamp 1623529830
transform 1 0 34500 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_372
timestamp 1623529830
transform 1 0 35328 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_384
timestamp 1623529830
transform 1 0 36432 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1623529830
transform -1 0 38824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_396
timestamp 1623529830
transform 1 0 37536 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_404
timestamp 1623529830
transform 1 0 38272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1623529830
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1623529830
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1623529830
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1623529830
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1623529830
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1623529830
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_51
timestamp 1623529830
transform 1 0 5796 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_58
timestamp 1623529830
transform 1 0 6440 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_70
timestamp 1623529830
transform 1 0 7544 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_82
timestamp 1623529830
transform 1 0 8648 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_94
timestamp 1623529830
transform 1 0 9752 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_106
timestamp 1623529830
transform 1 0 10856 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1623529830
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_115
timestamp 1623529830
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_127
timestamp 1623529830
transform 1 0 12788 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_139
timestamp 1623529830
transform 1 0 13892 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_151
timestamp 1623529830
transform 1 0 14996 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1623529830
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_163
timestamp 1623529830
transform 1 0 16100 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_172
timestamp 1623529830
transform 1 0 16928 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1623529830
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1623529830
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1623529830
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1623529830
transform 1 0 22080 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_220
timestamp 1623529830
transform 1 0 21344 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_229
timestamp 1623529830
transform 1 0 22172 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_241
timestamp 1623529830
transform 1 0 23276 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_253
timestamp 1623529830
transform 1 0 24380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_265
timestamp 1623529830
transform 1 0 25484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_277
timestamp 1623529830
transform 1 0 26588 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1623529830
transform 1 0 27324 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_286
timestamp 1623529830
transform 1 0 27416 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_298
timestamp 1623529830
transform 1 0 28520 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_310
timestamp 1623529830
transform 1 0 29624 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_322
timestamp 1623529830
transform 1 0 30728 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1623529830
transform 1 0 32568 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_334
timestamp 1623529830
transform 1 0 31832 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_343
timestamp 1623529830
transform 1 0 32660 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_355
timestamp 1623529830
transform 1 0 33764 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_367
timestamp 1623529830
transform 1 0 34868 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_379
timestamp 1623529830
transform 1 0 35972 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_391
timestamp 1623529830
transform 1 0 37076 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1623529830
transform -1 0 38824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1623529830
transform 1 0 37812 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_400
timestamp 1623529830
transform 1 0 37904 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_406
timestamp 1623529830
transform 1 0 38456 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1623529830
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1623529830
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1623529830
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1623529830
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1623529830
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_30
timestamp 1623529830
transform 1 0 3864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_42
timestamp 1623529830
transform 1 0 4968 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_54
timestamp 1623529830
transform 1 0 6072 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1623529830
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_66
timestamp 1623529830
transform 1 0 7176 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_78
timestamp 1623529830
transform 1 0 8280 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_87
timestamp 1623529830
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_99
timestamp 1623529830
transform 1 0 10212 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_111
timestamp 1623529830
transform 1 0 11316 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1623529830
transform 1 0 12420 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1623529830
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_135
timestamp 1623529830
transform 1 0 13524 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_144
timestamp 1623529830
transform 1 0 14352 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_156
timestamp 1623529830
transform 1 0 15456 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_168
timestamp 1623529830
transform 1 0 16560 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_180
timestamp 1623529830
transform 1 0 17664 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_192
timestamp 1623529830
transform 1 0 18768 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1623529830
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_201
timestamp 1623529830
transform 1 0 19596 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_213
timestamp 1623529830
transform 1 0 20700 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_225
timestamp 1623529830
transform 1 0 21804 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_237
timestamp 1623529830
transform 1 0 22908 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1623529830
transform 1 0 24748 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_249
timestamp 1623529830
transform 1 0 24012 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_258
timestamp 1623529830
transform 1 0 24840 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_270
timestamp 1623529830
transform 1 0 25944 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_282
timestamp 1623529830
transform 1 0 27048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_294
timestamp 1623529830
transform 1 0 28152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1623529830
transform 1 0 29992 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_306
timestamp 1623529830
transform 1 0 29256 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_315
timestamp 1623529830
transform 1 0 30084 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_327
timestamp 1623529830
transform 1 0 31188 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_339
timestamp 1623529830
transform 1 0 32292 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1623529830
transform 1 0 35236 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_351
timestamp 1623529830
transform 1 0 33396 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_363
timestamp 1623529830
transform 1 0 34500 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_372
timestamp 1623529830
transform 1 0 35328 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_384
timestamp 1623529830
transform 1 0 36432 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1623529830
transform -1 0 38824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_396
timestamp 1623529830
transform 1 0 37536 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_404
timestamp 1623529830
transform 1 0 38272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1623529830
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1623529830
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1623529830
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1623529830
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1623529830
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1623529830
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_51
timestamp 1623529830
transform 1 0 5796 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_58
timestamp 1623529830
transform 1 0 6440 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_70
timestamp 1623529830
transform 1 0 7544 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_82
timestamp 1623529830
transform 1 0 8648 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_94
timestamp 1623529830
transform 1 0 9752 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_106
timestamp 1623529830
transform 1 0 10856 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1623529830
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_115
timestamp 1623529830
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_127
timestamp 1623529830
transform 1 0 12788 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_139
timestamp 1623529830
transform 1 0 13892 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_151
timestamp 1623529830
transform 1 0 14996 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1623529830
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_163
timestamp 1623529830
transform 1 0 16100 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_172
timestamp 1623529830
transform 1 0 16928 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1623529830
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1623529830
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1623529830
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1623529830
transform 1 0 22080 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_220
timestamp 1623529830
transform 1 0 21344 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_229
timestamp 1623529830
transform 1 0 22172 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_241
timestamp 1623529830
transform 1 0 23276 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_253
timestamp 1623529830
transform 1 0 24380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_265
timestamp 1623529830
transform 1 0 25484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_277
timestamp 1623529830
transform 1 0 26588 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1623529830
transform 1 0 27324 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_286
timestamp 1623529830
transform 1 0 27416 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_298
timestamp 1623529830
transform 1 0 28520 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_310
timestamp 1623529830
transform 1 0 29624 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_322
timestamp 1623529830
transform 1 0 30728 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1623529830
transform 1 0 32568 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_334
timestamp 1623529830
transform 1 0 31832 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_343
timestamp 1623529830
transform 1 0 32660 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_355
timestamp 1623529830
transform 1 0 33764 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_367
timestamp 1623529830
transform 1 0 34868 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_379
timestamp 1623529830
transform 1 0 35972 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_391
timestamp 1623529830
transform 1 0 37076 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1623529830
transform -1 0 38824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1623529830
transform 1 0 37812 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_400
timestamp 1623529830
transform 1 0 37904 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_406
timestamp 1623529830
transform 1 0 38456 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1623529830
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1623529830
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1623529830
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1623529830
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1623529830
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1623529830
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1623529830
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1623529830
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_30
timestamp 1623529830
transform 1 0 3864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_42
timestamp 1623529830
transform 1 0 4968 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1623529830
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1623529830
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1623529830
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_54
timestamp 1623529830
transform 1 0 6072 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_51
timestamp 1623529830
transform 1 0 5796 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_58
timestamp 1623529830
transform 1 0 6440 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1623529830
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_66
timestamp 1623529830
transform 1 0 7176 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_78
timestamp 1623529830
transform 1 0 8280 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_87
timestamp 1623529830
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_70
timestamp 1623529830
transform 1 0 7544 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_82
timestamp 1623529830
transform 1 0 8648 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_99
timestamp 1623529830
transform 1 0 10212 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_94
timestamp 1623529830
transform 1 0 9752 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_106
timestamp 1623529830
transform 1 0 10856 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1623529830
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_111
timestamp 1623529830
transform 1 0 11316 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_123
timestamp 1623529830
transform 1 0 12420 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_115
timestamp 1623529830
transform 1 0 11684 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_127
timestamp 1623529830
transform 1 0 12788 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1623529830
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_135
timestamp 1623529830
transform 1 0 13524 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_144
timestamp 1623529830
transform 1 0 14352 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_139
timestamp 1623529830
transform 1 0 13892 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_151
timestamp 1623529830
transform 1 0 14996 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1623529830
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_156
timestamp 1623529830
transform 1 0 15456 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_168
timestamp 1623529830
transform 1 0 16560 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_163
timestamp 1623529830
transform 1 0 16100 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_172
timestamp 1623529830
transform 1 0 16928 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_180
timestamp 1623529830
transform 1 0 17664 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_192
timestamp 1623529830
transform 1 0 18768 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1623529830
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1623529830
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1623529830
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_201
timestamp 1623529830
transform 1 0 19596 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_213
timestamp 1623529830
transform 1 0 20700 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1623529830
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1623529830
transform 1 0 22080 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_225
timestamp 1623529830
transform 1 0 21804 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_237
timestamp 1623529830
transform 1 0 22908 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_220
timestamp 1623529830
transform 1 0 21344 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_229
timestamp 1623529830
transform 1 0 22172 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1623529830
transform 1 0 24748 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_249
timestamp 1623529830
transform 1 0 24012 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_258
timestamp 1623529830
transform 1 0 24840 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_241
timestamp 1623529830
transform 1 0 23276 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_253
timestamp 1623529830
transform 1 0 24380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_270
timestamp 1623529830
transform 1 0 25944 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_282
timestamp 1623529830
transform 1 0 27048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_265
timestamp 1623529830
transform 1 0 25484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_277
timestamp 1623529830
transform 1 0 26588 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1623529830
transform 1 0 27324 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_294
timestamp 1623529830
transform 1 0 28152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_286
timestamp 1623529830
transform 1 0 27416 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_298
timestamp 1623529830
transform 1 0 28520 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1623529830
transform 1 0 29992 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_306
timestamp 1623529830
transform 1 0 29256 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_315
timestamp 1623529830
transform 1 0 30084 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_327
timestamp 1623529830
transform 1 0 31188 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_310
timestamp 1623529830
transform 1 0 29624 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_322
timestamp 1623529830
transform 1 0 30728 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1623529830
transform 1 0 32568 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_339
timestamp 1623529830
transform 1 0 32292 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_334
timestamp 1623529830
transform 1 0 31832 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_343
timestamp 1623529830
transform 1 0 32660 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1623529830
transform 1 0 35236 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_351
timestamp 1623529830
transform 1 0 33396 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_363
timestamp 1623529830
transform 1 0 34500 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_355
timestamp 1623529830
transform 1 0 33764 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_367
timestamp 1623529830
transform 1 0 34868 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_372
timestamp 1623529830
transform 1 0 35328 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_384
timestamp 1623529830
transform 1 0 36432 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_379
timestamp 1623529830
transform 1 0 35972 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_391
timestamp 1623529830
transform 1 0 37076 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1623529830
transform -1 0 38824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1623529830
transform -1 0 38824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1623529830
transform 1 0 37812 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_396
timestamp 1623529830
transform 1 0 37536 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_404
timestamp 1623529830
transform 1 0 38272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_400
timestamp 1623529830
transform 1 0 37904 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_406
timestamp 1623529830
transform 1 0 38456 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1623529830
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1623529830
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1623529830
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1623529830
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1623529830
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_30
timestamp 1623529830
transform 1 0 3864 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_42
timestamp 1623529830
transform 1 0 4968 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_54
timestamp 1623529830
transform 1 0 6072 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1623529830
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_66
timestamp 1623529830
transform 1 0 7176 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_78
timestamp 1623529830
transform 1 0 8280 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_87
timestamp 1623529830
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_99
timestamp 1623529830
transform 1 0 10212 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_111
timestamp 1623529830
transform 1 0 11316 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_123
timestamp 1623529830
transform 1 0 12420 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1623529830
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_135
timestamp 1623529830
transform 1 0 13524 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_144
timestamp 1623529830
transform 1 0 14352 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_156
timestamp 1623529830
transform 1 0 15456 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_168
timestamp 1623529830
transform 1 0 16560 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_180
timestamp 1623529830
transform 1 0 17664 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_192
timestamp 1623529830
transform 1 0 18768 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1623529830
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_201
timestamp 1623529830
transform 1 0 19596 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_213
timestamp 1623529830
transform 1 0 20700 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_225
timestamp 1623529830
transform 1 0 21804 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_237
timestamp 1623529830
transform 1 0 22908 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1623529830
transform 1 0 24748 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_249
timestamp 1623529830
transform 1 0 24012 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_258
timestamp 1623529830
transform 1 0 24840 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_270
timestamp 1623529830
transform 1 0 25944 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_282
timestamp 1623529830
transform 1 0 27048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_294
timestamp 1623529830
transform 1 0 28152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1623529830
transform 1 0 29992 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_306
timestamp 1623529830
transform 1 0 29256 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_315
timestamp 1623529830
transform 1 0 30084 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_327
timestamp 1623529830
transform 1 0 31188 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_339
timestamp 1623529830
transform 1 0 32292 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1623529830
transform 1 0 35236 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_351
timestamp 1623529830
transform 1 0 33396 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_363
timestamp 1623529830
transform 1 0 34500 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_372
timestamp 1623529830
transform 1 0 35328 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_384
timestamp 1623529830
transform 1 0 36432 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1623529830
transform -1 0 38824 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_396
timestamp 1623529830
transform 1 0 37536 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_404
timestamp 1623529830
transform 1 0 38272 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1623529830
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1623529830
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1623529830
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1623529830
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1623529830
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1623529830
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_51
timestamp 1623529830
transform 1 0 5796 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_58
timestamp 1623529830
transform 1 0 6440 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_70
timestamp 1623529830
transform 1 0 7544 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_82
timestamp 1623529830
transform 1 0 8648 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_94
timestamp 1623529830
transform 1 0 9752 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_106
timestamp 1623529830
transform 1 0 10856 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1623529830
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_115
timestamp 1623529830
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_127
timestamp 1623529830
transform 1 0 12788 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_139
timestamp 1623529830
transform 1 0 13892 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_151
timestamp 1623529830
transform 1 0 14996 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1623529830
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_163
timestamp 1623529830
transform 1 0 16100 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_172
timestamp 1623529830
transform 1 0 16928 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1623529830
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1623529830
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1623529830
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1623529830
transform 1 0 22080 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_220
timestamp 1623529830
transform 1 0 21344 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_229
timestamp 1623529830
transform 1 0 22172 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_241
timestamp 1623529830
transform 1 0 23276 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_253
timestamp 1623529830
transform 1 0 24380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_265
timestamp 1623529830
transform 1 0 25484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_277
timestamp 1623529830
transform 1 0 26588 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1623529830
transform 1 0 27324 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_286
timestamp 1623529830
transform 1 0 27416 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_298
timestamp 1623529830
transform 1 0 28520 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_310
timestamp 1623529830
transform 1 0 29624 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_322
timestamp 1623529830
transform 1 0 30728 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1623529830
transform 1 0 32568 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_334
timestamp 1623529830
transform 1 0 31832 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_343
timestamp 1623529830
transform 1 0 32660 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_355
timestamp 1623529830
transform 1 0 33764 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_367
timestamp 1623529830
transform 1 0 34868 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_379
timestamp 1623529830
transform 1 0 35972 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_391
timestamp 1623529830
transform 1 0 37076 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1623529830
transform -1 0 38824 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1623529830
transform 1 0 37812 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_400
timestamp 1623529830
transform 1 0 37904 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_406
timestamp 1623529830
transform 1 0 38456 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1623529830
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1623529830
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1623529830
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1623529830
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1623529830
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_30
timestamp 1623529830
transform 1 0 3864 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_42
timestamp 1623529830
transform 1 0 4968 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_54
timestamp 1623529830
transform 1 0 6072 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1623529830
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_66
timestamp 1623529830
transform 1 0 7176 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_78
timestamp 1623529830
transform 1 0 8280 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_87
timestamp 1623529830
transform 1 0 9108 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_99
timestamp 1623529830
transform 1 0 10212 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_111
timestamp 1623529830
transform 1 0 11316 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_123
timestamp 1623529830
transform 1 0 12420 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1623529830
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_135
timestamp 1623529830
transform 1 0 13524 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_144
timestamp 1623529830
transform 1 0 14352 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_156
timestamp 1623529830
transform 1 0 15456 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_168
timestamp 1623529830
transform 1 0 16560 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_180
timestamp 1623529830
transform 1 0 17664 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_192
timestamp 1623529830
transform 1 0 18768 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1623529830
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_201
timestamp 1623529830
transform 1 0 19596 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_213
timestamp 1623529830
transform 1 0 20700 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_225
timestamp 1623529830
transform 1 0 21804 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_237
timestamp 1623529830
transform 1 0 22908 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1623529830
transform 1 0 24748 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_249
timestamp 1623529830
transform 1 0 24012 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_258
timestamp 1623529830
transform 1 0 24840 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_270
timestamp 1623529830
transform 1 0 25944 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_282
timestamp 1623529830
transform 1 0 27048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_294
timestamp 1623529830
transform 1 0 28152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1623529830
transform 1 0 29992 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_306
timestamp 1623529830
transform 1 0 29256 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_315
timestamp 1623529830
transform 1 0 30084 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_327
timestamp 1623529830
transform 1 0 31188 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_339
timestamp 1623529830
transform 1 0 32292 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1623529830
transform 1 0 35236 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_351
timestamp 1623529830
transform 1 0 33396 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_363
timestamp 1623529830
transform 1 0 34500 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_372
timestamp 1623529830
transform 1 0 35328 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_384
timestamp 1623529830
transform 1 0 36432 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1623529830
transform -1 0 38824 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_396
timestamp 1623529830
transform 1 0 37536 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_404
timestamp 1623529830
transform 1 0 38272 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1623529830
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1623529830
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1623529830
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1623529830
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1623529830
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1623529830
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_51
timestamp 1623529830
transform 1 0 5796 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_58
timestamp 1623529830
transform 1 0 6440 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_70
timestamp 1623529830
transform 1 0 7544 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_82
timestamp 1623529830
transform 1 0 8648 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_94
timestamp 1623529830
transform 1 0 9752 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_106
timestamp 1623529830
transform 1 0 10856 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1623529830
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_115
timestamp 1623529830
transform 1 0 11684 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_127
timestamp 1623529830
transform 1 0 12788 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_139
timestamp 1623529830
transform 1 0 13892 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_151
timestamp 1623529830
transform 1 0 14996 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1623529830
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_163
timestamp 1623529830
transform 1 0 16100 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_172
timestamp 1623529830
transform 1 0 16928 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1623529830
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1623529830
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1623529830
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1623529830
transform 1 0 22080 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_220
timestamp 1623529830
transform 1 0 21344 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_229
timestamp 1623529830
transform 1 0 22172 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_241
timestamp 1623529830
transform 1 0 23276 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_253
timestamp 1623529830
transform 1 0 24380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_265
timestamp 1623529830
transform 1 0 25484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_277
timestamp 1623529830
transform 1 0 26588 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1623529830
transform 1 0 27324 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_286
timestamp 1623529830
transform 1 0 27416 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_298
timestamp 1623529830
transform 1 0 28520 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_310
timestamp 1623529830
transform 1 0 29624 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_322
timestamp 1623529830
transform 1 0 30728 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1623529830
transform 1 0 32568 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_334
timestamp 1623529830
transform 1 0 31832 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_343
timestamp 1623529830
transform 1 0 32660 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_355
timestamp 1623529830
transform 1 0 33764 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_367
timestamp 1623529830
transform 1 0 34868 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_379
timestamp 1623529830
transform 1 0 35972 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_391
timestamp 1623529830
transform 1 0 37076 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1623529830
transform -1 0 38824 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1623529830
transform 1 0 37812 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_400
timestamp 1623529830
transform 1 0 37904 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_406
timestamp 1623529830
transform 1 0 38456 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1623529830
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1623529830
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1623529830
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1623529830
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_27
timestamp 1623529830
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_30
timestamp 1623529830
transform 1 0 3864 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_42
timestamp 1623529830
transform 1 0 4968 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_54
timestamp 1623529830
transform 1 0 6072 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1623529830
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_66
timestamp 1623529830
transform 1 0 7176 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_78
timestamp 1623529830
transform 1 0 8280 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_87
timestamp 1623529830
transform 1 0 9108 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_99
timestamp 1623529830
transform 1 0 10212 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_111
timestamp 1623529830
transform 1 0 11316 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_123
timestamp 1623529830
transform 1 0 12420 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1623529830
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_135
timestamp 1623529830
transform 1 0 13524 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_144
timestamp 1623529830
transform 1 0 14352 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1623529830
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1623529830
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_180
timestamp 1623529830
transform 1 0 17664 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_192
timestamp 1623529830
transform 1 0 18768 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1623529830
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_201
timestamp 1623529830
transform 1 0 19596 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_213
timestamp 1623529830
transform 1 0 20700 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_225
timestamp 1623529830
transform 1 0 21804 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_237
timestamp 1623529830
transform 1 0 22908 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1623529830
transform 1 0 24748 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_249
timestamp 1623529830
transform 1 0 24012 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_258
timestamp 1623529830
transform 1 0 24840 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_270
timestamp 1623529830
transform 1 0 25944 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_282
timestamp 1623529830
transform 1 0 27048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_294
timestamp 1623529830
transform 1 0 28152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1623529830
transform 1 0 29992 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_306
timestamp 1623529830
transform 1 0 29256 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_315
timestamp 1623529830
transform 1 0 30084 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_327
timestamp 1623529830
transform 1 0 31188 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_339
timestamp 1623529830
transform 1 0 32292 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1623529830
transform 1 0 35236 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_351
timestamp 1623529830
transform 1 0 33396 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_363
timestamp 1623529830
transform 1 0 34500 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_372
timestamp 1623529830
transform 1 0 35328 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_384
timestamp 1623529830
transform 1 0 36432 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1623529830
transform -1 0 38824 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623529830
transform -1 0 38180 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_396
timestamp 1623529830
transform 1 0 37536 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_403
timestamp 1623529830
transform 1 0 38180 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1623529830
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1623529830
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1623529830
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1623529830
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1623529830
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1623529830
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1623529830
transform 1 0 3772 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1623529830
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1623529830
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1623529830
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_30
timestamp 1623529830
transform 1 0 3864 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_42
timestamp 1623529830
transform 1 0 4968 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1623529830
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_51
timestamp 1623529830
transform 1 0 5796 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_58
timestamp 1623529830
transform 1 0 6440 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_54
timestamp 1623529830
transform 1 0 6072 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1623529830
transform 1 0 9016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_70
timestamp 1623529830
transform 1 0 7544 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_82
timestamp 1623529830
transform 1 0 8648 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_66
timestamp 1623529830
transform 1 0 7176 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_78
timestamp 1623529830
transform 1 0 8280 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_87
timestamp 1623529830
transform 1 0 9108 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_94
timestamp 1623529830
transform 1 0 9752 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_106
timestamp 1623529830
transform 1 0 10856 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_99
timestamp 1623529830
transform 1 0 10212 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1623529830
transform 1 0 11592 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_115
timestamp 1623529830
transform 1 0 11684 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_127
timestamp 1623529830
transform 1 0 12788 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_111
timestamp 1623529830
transform 1 0 11316 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_123
timestamp 1623529830
transform 1 0 12420 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1623529830
transform 1 0 14260 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_139
timestamp 1623529830
transform 1 0 13892 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_151
timestamp 1623529830
transform 1 0 14996 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_135
timestamp 1623529830
transform 1 0 13524 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_144
timestamp 1623529830
transform 1 0 14352 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1623529830
transform 1 0 16836 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_163
timestamp 1623529830
transform 1 0 16100 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_172
timestamp 1623529830
transform 1 0 16928 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_156
timestamp 1623529830
transform 1 0 15456 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_168
timestamp 1623529830
transform 1 0 16560 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1623529830
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1623529830
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_180
timestamp 1623529830
transform 1 0 17664 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_192
timestamp 1623529830
transform 1 0 18768 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1623529830
transform 1 0 19504 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1623529830
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_201
timestamp 1623529830
transform 1 0 19596 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_213
timestamp 1623529830
transform 1 0 20700 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1623529830
transform 1 0 22080 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_220
timestamp 1623529830
transform 1 0 21344 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_229
timestamp 1623529830
transform 1 0 22172 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_225
timestamp 1623529830
transform 1 0 21804 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_237
timestamp 1623529830
transform 1 0 22908 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1623529830
transform 1 0 24748 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_241
timestamp 1623529830
transform 1 0 23276 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_253
timestamp 1623529830
transform 1 0 24380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_249
timestamp 1623529830
transform 1 0 24012 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_258
timestamp 1623529830
transform 1 0 24840 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_265
timestamp 1623529830
transform 1 0 25484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_277
timestamp 1623529830
transform 1 0 26588 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_270
timestamp 1623529830
transform 1 0 25944 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_282
timestamp 1623529830
transform 1 0 27048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1623529830
transform 1 0 27324 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_286
timestamp 1623529830
transform 1 0 27416 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_298
timestamp 1623529830
transform 1 0 28520 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_294
timestamp 1623529830
transform 1 0 28152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1623529830
transform 1 0 29992 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_310
timestamp 1623529830
transform 1 0 29624 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_322
timestamp 1623529830
transform 1 0 30728 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_306
timestamp 1623529830
transform 1 0 29256 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_315
timestamp 1623529830
transform 1 0 30084 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_327
timestamp 1623529830
transform 1 0 31188 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1623529830
transform 1 0 32568 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_334
timestamp 1623529830
transform 1 0 31832 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_343
timestamp 1623529830
transform 1 0 32660 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_339
timestamp 1623529830
transform 1 0 32292 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1623529830
transform 1 0 35236 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_355
timestamp 1623529830
transform 1 0 33764 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_367
timestamp 1623529830
transform 1 0 34868 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_351
timestamp 1623529830
transform 1 0 33396 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_363
timestamp 1623529830
transform 1 0 34500 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_379
timestamp 1623529830
transform 1 0 35972 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_391
timestamp 1623529830
transform 1 0 37076 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_372
timestamp 1623529830
transform 1 0 35328 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_384
timestamp 1623529830
transform 1 0 36432 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1623529830
transform -1 0 38824 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1623529830
transform -1 0 38824 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1623529830
transform 1 0 37812 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_400
timestamp 1623529830
transform 1 0 37904 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_406
timestamp 1623529830
transform 1 0 38456 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_396
timestamp 1623529830
transform 1 0 37536 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_404
timestamp 1623529830
transform 1 0 38272 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1623529830
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1623529830
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1623529830
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1623529830
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1623529830
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1623529830
transform 1 0 6348 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_51
timestamp 1623529830
transform 1 0 5796 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_58
timestamp 1623529830
transform 1 0 6440 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_70
timestamp 1623529830
transform 1 0 7544 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_82
timestamp 1623529830
transform 1 0 8648 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1623529830
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_106
timestamp 1623529830
transform 1 0 10856 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1623529830
transform 1 0 11592 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_115
timestamp 1623529830
transform 1 0 11684 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_127
timestamp 1623529830
transform 1 0 12788 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_139
timestamp 1623529830
transform 1 0 13892 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_151
timestamp 1623529830
transform 1 0 14996 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1623529830
transform 1 0 16836 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_163
timestamp 1623529830
transform 1 0 16100 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_172
timestamp 1623529830
transform 1 0 16928 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1623529830
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1623529830
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1623529830
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1623529830
transform 1 0 22080 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_220
timestamp 1623529830
transform 1 0 21344 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_229
timestamp 1623529830
transform 1 0 22172 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_241
timestamp 1623529830
transform 1 0 23276 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_253
timestamp 1623529830
transform 1 0 24380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_265
timestamp 1623529830
transform 1 0 25484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_277
timestamp 1623529830
transform 1 0 26588 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1623529830
transform 1 0 27324 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_286
timestamp 1623529830
transform 1 0 27416 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_298
timestamp 1623529830
transform 1 0 28520 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_310
timestamp 1623529830
transform 1 0 29624 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_322
timestamp 1623529830
transform 1 0 30728 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1623529830
transform 1 0 32568 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_334
timestamp 1623529830
transform 1 0 31832 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_343
timestamp 1623529830
transform 1 0 32660 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_355
timestamp 1623529830
transform 1 0 33764 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_367
timestamp 1623529830
transform 1 0 34868 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_379
timestamp 1623529830
transform 1 0 35972 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_391
timestamp 1623529830
transform 1 0 37076 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1623529830
transform -1 0 38824 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1623529830
transform 1 0 37812 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_400
timestamp 1623529830
transform 1 0 37904 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_406
timestamp 1623529830
transform 1 0 38456 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1623529830
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1623529830
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1623529830
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1623529830
transform 1 0 3772 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1623529830
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_30
timestamp 1623529830
transform 1 0 3864 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_42
timestamp 1623529830
transform 1 0 4968 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_54
timestamp 1623529830
transform 1 0 6072 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1623529830
transform 1 0 9016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_66
timestamp 1623529830
transform 1 0 7176 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_78
timestamp 1623529830
transform 1 0 8280 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_87
timestamp 1623529830
transform 1 0 9108 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_99
timestamp 1623529830
transform 1 0 10212 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_111
timestamp 1623529830
transform 1 0 11316 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_123
timestamp 1623529830
transform 1 0 12420 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1623529830
transform 1 0 14260 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_135
timestamp 1623529830
transform 1 0 13524 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_144
timestamp 1623529830
transform 1 0 14352 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_156
timestamp 1623529830
transform 1 0 15456 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_168
timestamp 1623529830
transform 1 0 16560 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_180
timestamp 1623529830
transform 1 0 17664 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_192
timestamp 1623529830
transform 1 0 18768 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1623529830
transform 1 0 19504 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_201
timestamp 1623529830
transform 1 0 19596 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_213
timestamp 1623529830
transform 1 0 20700 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_225
timestamp 1623529830
transform 1 0 21804 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_237
timestamp 1623529830
transform 1 0 22908 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1623529830
transform 1 0 24748 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_249
timestamp 1623529830
transform 1 0 24012 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_258
timestamp 1623529830
transform 1 0 24840 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_270
timestamp 1623529830
transform 1 0 25944 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_282
timestamp 1623529830
transform 1 0 27048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_294
timestamp 1623529830
transform 1 0 28152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1623529830
transform 1 0 29992 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_306
timestamp 1623529830
transform 1 0 29256 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_315
timestamp 1623529830
transform 1 0 30084 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_327
timestamp 1623529830
transform 1 0 31188 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_339
timestamp 1623529830
transform 1 0 32292 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1623529830
transform 1 0 35236 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_351
timestamp 1623529830
transform 1 0 33396 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_363
timestamp 1623529830
transform 1 0 34500 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_372
timestamp 1623529830
transform 1 0 35328 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_384
timestamp 1623529830
transform 1 0 36432 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1623529830
transform -1 0 38824 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_396
timestamp 1623529830
transform 1 0 37536 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_404
timestamp 1623529830
transform 1 0 38272 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1623529830
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1623529830
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1623529830
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1623529830
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1623529830
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1623529830
transform 1 0 6348 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_51
timestamp 1623529830
transform 1 0 5796 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_58
timestamp 1623529830
transform 1 0 6440 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_70
timestamp 1623529830
transform 1 0 7544 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_82
timestamp 1623529830
transform 1 0 8648 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_94
timestamp 1623529830
transform 1 0 9752 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_106
timestamp 1623529830
transform 1 0 10856 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1623529830
transform 1 0 11592 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_115
timestamp 1623529830
transform 1 0 11684 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_127
timestamp 1623529830
transform 1 0 12788 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_139
timestamp 1623529830
transform 1 0 13892 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_151
timestamp 1623529830
transform 1 0 14996 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1623529830
transform 1 0 16836 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_163
timestamp 1623529830
transform 1 0 16100 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_172
timestamp 1623529830
transform 1 0 16928 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1623529830
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1623529830
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1623529830
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1623529830
transform 1 0 22080 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_220
timestamp 1623529830
transform 1 0 21344 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_229
timestamp 1623529830
transform 1 0 22172 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_241
timestamp 1623529830
transform 1 0 23276 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_253
timestamp 1623529830
transform 1 0 24380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_265
timestamp 1623529830
transform 1 0 25484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_277
timestamp 1623529830
transform 1 0 26588 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1623529830
transform 1 0 27324 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_286
timestamp 1623529830
transform 1 0 27416 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_298
timestamp 1623529830
transform 1 0 28520 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_310
timestamp 1623529830
transform 1 0 29624 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_322
timestamp 1623529830
transform 1 0 30728 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1623529830
transform 1 0 32568 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_334
timestamp 1623529830
transform 1 0 31832 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_343
timestamp 1623529830
transform 1 0 32660 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_355
timestamp 1623529830
transform 1 0 33764 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_367
timestamp 1623529830
transform 1 0 34868 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_379
timestamp 1623529830
transform 1 0 35972 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_391
timestamp 1623529830
transform 1 0 37076 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1623529830
transform -1 0 38824 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1623529830
transform 1 0 37812 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_400
timestamp 1623529830
transform 1 0 37904 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_406
timestamp 1623529830
transform 1 0 38456 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1623529830
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1623529830
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1623529830
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1623529830
transform 1 0 3772 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_27
timestamp 1623529830
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_30
timestamp 1623529830
transform 1 0 3864 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_42
timestamp 1623529830
transform 1 0 4968 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_54
timestamp 1623529830
transform 1 0 6072 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1623529830
transform 1 0 9016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_66
timestamp 1623529830
transform 1 0 7176 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_78
timestamp 1623529830
transform 1 0 8280 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_87
timestamp 1623529830
transform 1 0 9108 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_99
timestamp 1623529830
transform 1 0 10212 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_111
timestamp 1623529830
transform 1 0 11316 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_123
timestamp 1623529830
transform 1 0 12420 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1623529830
transform 1 0 14260 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_135
timestamp 1623529830
transform 1 0 13524 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_144
timestamp 1623529830
transform 1 0 14352 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_156
timestamp 1623529830
transform 1 0 15456 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_168
timestamp 1623529830
transform 1 0 16560 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_180
timestamp 1623529830
transform 1 0 17664 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_192
timestamp 1623529830
transform 1 0 18768 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1623529830
transform 1 0 19504 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_201
timestamp 1623529830
transform 1 0 19596 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_213
timestamp 1623529830
transform 1 0 20700 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_225
timestamp 1623529830
transform 1 0 21804 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_237
timestamp 1623529830
transform 1 0 22908 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1623529830
transform 1 0 24748 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_249
timestamp 1623529830
transform 1 0 24012 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_258
timestamp 1623529830
transform 1 0 24840 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_270
timestamp 1623529830
transform 1 0 25944 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_282
timestamp 1623529830
transform 1 0 27048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_294
timestamp 1623529830
transform 1 0 28152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1623529830
transform 1 0 29992 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_306
timestamp 1623529830
transform 1 0 29256 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_315
timestamp 1623529830
transform 1 0 30084 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_327
timestamp 1623529830
transform 1 0 31188 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_339
timestamp 1623529830
transform 1 0 32292 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1623529830
transform 1 0 35236 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_351
timestamp 1623529830
transform 1 0 33396 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_363
timestamp 1623529830
transform 1 0 34500 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_372
timestamp 1623529830
transform 1 0 35328 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_384
timestamp 1623529830
transform 1 0 36432 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1623529830
transform -1 0 38824 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_396
timestamp 1623529830
transform 1 0 37536 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_404
timestamp 1623529830
transform 1 0 38272 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1623529830
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1623529830
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1623529830
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1623529830
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1623529830
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1623529830
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1623529830
transform 1 0 3772 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1623529830
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1623529830
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_27
timestamp 1623529830
transform 1 0 3588 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_30
timestamp 1623529830
transform 1 0 3864 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_42
timestamp 1623529830
transform 1 0 4968 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1623529830
transform 1 0 6348 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_51
timestamp 1623529830
transform 1 0 5796 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_58
timestamp 1623529830
transform 1 0 6440 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_54
timestamp 1623529830
transform 1 0 6072 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1623529830
transform 1 0 9016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_70
timestamp 1623529830
transform 1 0 7544 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_82
timestamp 1623529830
transform 1 0 8648 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_66
timestamp 1623529830
transform 1 0 7176 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_78
timestamp 1623529830
transform 1 0 8280 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_87
timestamp 1623529830
transform 1 0 9108 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_94
timestamp 1623529830
transform 1 0 9752 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_106
timestamp 1623529830
transform 1 0 10856 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_99
timestamp 1623529830
transform 1 0 10212 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1623529830
transform 1 0 11592 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_115
timestamp 1623529830
transform 1 0 11684 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_127
timestamp 1623529830
transform 1 0 12788 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_111
timestamp 1623529830
transform 1 0 11316 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_123
timestamp 1623529830
transform 1 0 12420 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1623529830
transform 1 0 14260 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_139
timestamp 1623529830
transform 1 0 13892 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_151
timestamp 1623529830
transform 1 0 14996 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_135
timestamp 1623529830
transform 1 0 13524 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_144
timestamp 1623529830
transform 1 0 14352 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1623529830
transform 1 0 16836 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_163
timestamp 1623529830
transform 1 0 16100 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_172
timestamp 1623529830
transform 1 0 16928 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_156
timestamp 1623529830
transform 1 0 15456 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_168
timestamp 1623529830
transform 1 0 16560 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1623529830
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_196
timestamp 1623529830
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_180
timestamp 1623529830
transform 1 0 17664 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_192
timestamp 1623529830
transform 1 0 18768 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1623529830
transform 1 0 19504 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1623529830
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_201
timestamp 1623529830
transform 1 0 19596 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_213
timestamp 1623529830
transform 1 0 20700 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1623529830
transform 1 0 22080 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_220
timestamp 1623529830
transform 1 0 21344 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_229
timestamp 1623529830
transform 1 0 22172 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_225
timestamp 1623529830
transform 1 0 21804 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_237
timestamp 1623529830
transform 1 0 22908 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1623529830
transform 1 0 24748 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_241
timestamp 1623529830
transform 1 0 23276 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_253
timestamp 1623529830
transform 1 0 24380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_249
timestamp 1623529830
transform 1 0 24012 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_258
timestamp 1623529830
transform 1 0 24840 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_265
timestamp 1623529830
transform 1 0 25484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_277
timestamp 1623529830
transform 1 0 26588 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_270
timestamp 1623529830
transform 1 0 25944 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_282
timestamp 1623529830
transform 1 0 27048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1623529830
transform 1 0 27324 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_286
timestamp 1623529830
transform 1 0 27416 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_298
timestamp 1623529830
transform 1 0 28520 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_294
timestamp 1623529830
transform 1 0 28152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1623529830
transform 1 0 29992 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_310
timestamp 1623529830
transform 1 0 29624 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_322
timestamp 1623529830
transform 1 0 30728 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_306
timestamp 1623529830
transform 1 0 29256 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_315
timestamp 1623529830
transform 1 0 30084 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_327
timestamp 1623529830
transform 1 0 31188 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1623529830
transform 1 0 32568 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_334
timestamp 1623529830
transform 1 0 31832 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_343
timestamp 1623529830
transform 1 0 32660 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_339
timestamp 1623529830
transform 1 0 32292 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1623529830
transform 1 0 35236 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_355
timestamp 1623529830
transform 1 0 33764 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_367
timestamp 1623529830
transform 1 0 34868 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_351
timestamp 1623529830
transform 1 0 33396 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_363
timestamp 1623529830
transform 1 0 34500 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_379
timestamp 1623529830
transform 1 0 35972 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_391
timestamp 1623529830
transform 1 0 37076 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_372
timestamp 1623529830
transform 1 0 35328 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_384
timestamp 1623529830
transform 1 0 36432 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1623529830
transform -1 0 38824 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1623529830
transform -1 0 38824 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1623529830
transform 1 0 37812 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_400
timestamp 1623529830
transform 1 0 37904 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_406
timestamp 1623529830
transform 1 0 38456 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_396
timestamp 1623529830
transform 1 0 37536 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_404
timestamp 1623529830
transform 1 0 38272 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1623529830
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1623529830
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1623529830
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1623529830
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1623529830
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1623529830
transform 1 0 6348 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_51
timestamp 1623529830
transform 1 0 5796 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_58
timestamp 1623529830
transform 1 0 6440 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_70
timestamp 1623529830
transform 1 0 7544 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_82
timestamp 1623529830
transform 1 0 8648 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_94
timestamp 1623529830
transform 1 0 9752 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_106
timestamp 1623529830
transform 1 0 10856 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1623529830
transform 1 0 11592 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_115
timestamp 1623529830
transform 1 0 11684 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_127
timestamp 1623529830
transform 1 0 12788 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_139
timestamp 1623529830
transform 1 0 13892 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_151
timestamp 1623529830
transform 1 0 14996 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1623529830
transform 1 0 16836 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_163
timestamp 1623529830
transform 1 0 16100 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_172
timestamp 1623529830
transform 1 0 16928 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1623529830
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1623529830
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1623529830
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1623529830
transform 1 0 22080 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_220
timestamp 1623529830
transform 1 0 21344 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_229
timestamp 1623529830
transform 1 0 22172 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_241
timestamp 1623529830
transform 1 0 23276 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_253
timestamp 1623529830
transform 1 0 24380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_265
timestamp 1623529830
transform 1 0 25484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_277
timestamp 1623529830
transform 1 0 26588 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1623529830
transform 1 0 27324 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_286
timestamp 1623529830
transform 1 0 27416 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_298
timestamp 1623529830
transform 1 0 28520 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_310
timestamp 1623529830
transform 1 0 29624 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_322
timestamp 1623529830
transform 1 0 30728 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1623529830
transform 1 0 32568 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_334
timestamp 1623529830
transform 1 0 31832 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_343
timestamp 1623529830
transform 1 0 32660 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_355
timestamp 1623529830
transform 1 0 33764 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_367
timestamp 1623529830
transform 1 0 34868 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_379
timestamp 1623529830
transform 1 0 35972 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_391
timestamp 1623529830
transform 1 0 37076 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1623529830
transform -1 0 38824 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1623529830
transform 1 0 37812 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_400
timestamp 1623529830
transform 1 0 37904 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_406
timestamp 1623529830
transform 1 0 38456 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1623529830
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1623529830
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1623529830
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1623529830
transform 1 0 3772 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_27
timestamp 1623529830
transform 1 0 3588 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_30
timestamp 1623529830
transform 1 0 3864 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_42
timestamp 1623529830
transform 1 0 4968 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_54
timestamp 1623529830
transform 1 0 6072 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1623529830
transform 1 0 9016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_66
timestamp 1623529830
transform 1 0 7176 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_78
timestamp 1623529830
transform 1 0 8280 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_87
timestamp 1623529830
transform 1 0 9108 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_99
timestamp 1623529830
transform 1 0 10212 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_111
timestamp 1623529830
transform 1 0 11316 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_123
timestamp 1623529830
transform 1 0 12420 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1623529830
transform 1 0 14260 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_135
timestamp 1623529830
transform 1 0 13524 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_144
timestamp 1623529830
transform 1 0 14352 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1623529830
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1623529830
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_180
timestamp 1623529830
transform 1 0 17664 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_192
timestamp 1623529830
transform 1 0 18768 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1623529830
transform 1 0 19504 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_201
timestamp 1623529830
transform 1 0 19596 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_213
timestamp 1623529830
transform 1 0 20700 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_225
timestamp 1623529830
transform 1 0 21804 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_237
timestamp 1623529830
transform 1 0 22908 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1623529830
transform 1 0 24748 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_249
timestamp 1623529830
transform 1 0 24012 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_258
timestamp 1623529830
transform 1 0 24840 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_270
timestamp 1623529830
transform 1 0 25944 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_282
timestamp 1623529830
transform 1 0 27048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_294
timestamp 1623529830
transform 1 0 28152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1623529830
transform 1 0 29992 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_306
timestamp 1623529830
transform 1 0 29256 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_315
timestamp 1623529830
transform 1 0 30084 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_327
timestamp 1623529830
transform 1 0 31188 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_339
timestamp 1623529830
transform 1 0 32292 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1623529830
transform 1 0 35236 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_351
timestamp 1623529830
transform 1 0 33396 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_363
timestamp 1623529830
transform 1 0 34500 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_372
timestamp 1623529830
transform 1 0 35328 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_384
timestamp 1623529830
transform 1 0 36432 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1623529830
transform -1 0 38824 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_396
timestamp 1623529830
transform 1 0 37536 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_404
timestamp 1623529830
transform 1 0 38272 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1623529830
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1623529830
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1623529830
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1623529830
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1623529830
transform 1 0 4692 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1623529830
transform 1 0 6348 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_51
timestamp 1623529830
transform 1 0 5796 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_58
timestamp 1623529830
transform 1 0 6440 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_70
timestamp 1623529830
transform 1 0 7544 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_82
timestamp 1623529830
transform 1 0 8648 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_94
timestamp 1623529830
transform 1 0 9752 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_106
timestamp 1623529830
transform 1 0 10856 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1623529830
transform 1 0 11592 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_115
timestamp 1623529830
transform 1 0 11684 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_127
timestamp 1623529830
transform 1 0 12788 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_139
timestamp 1623529830
transform 1 0 13892 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_151
timestamp 1623529830
transform 1 0 14996 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1623529830
transform 1 0 16836 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_163
timestamp 1623529830
transform 1 0 16100 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_172
timestamp 1623529830
transform 1 0 16928 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_184
timestamp 1623529830
transform 1 0 18032 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_196
timestamp 1623529830
transform 1 0 19136 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_208
timestamp 1623529830
transform 1 0 20240 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1623529830
transform 1 0 22080 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_220
timestamp 1623529830
transform 1 0 21344 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_229
timestamp 1623529830
transform 1 0 22172 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_241
timestamp 1623529830
transform 1 0 23276 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_253
timestamp 1623529830
transform 1 0 24380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_265
timestamp 1623529830
transform 1 0 25484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_277
timestamp 1623529830
transform 1 0 26588 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1623529830
transform 1 0 27324 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_286
timestamp 1623529830
transform 1 0 27416 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_298
timestamp 1623529830
transform 1 0 28520 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_310
timestamp 1623529830
transform 1 0 29624 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_322
timestamp 1623529830
transform 1 0 30728 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1623529830
transform 1 0 32568 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_334
timestamp 1623529830
transform 1 0 31832 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_343
timestamp 1623529830
transform 1 0 32660 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_355
timestamp 1623529830
transform 1 0 33764 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_367
timestamp 1623529830
transform 1 0 34868 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_379
timestamp 1623529830
transform 1 0 35972 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_391
timestamp 1623529830
transform 1 0 37076 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1623529830
transform -1 0 38824 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1623529830
transform 1 0 37812 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_400
timestamp 1623529830
transform 1 0 37904 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_406
timestamp 1623529830
transform 1 0 38456 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1623529830
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1623529830
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1623529830
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1623529830
transform 1 0 3772 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_27
timestamp 1623529830
transform 1 0 3588 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_30
timestamp 1623529830
transform 1 0 3864 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_42
timestamp 1623529830
transform 1 0 4968 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_54
timestamp 1623529830
transform 1 0 6072 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1623529830
transform 1 0 9016 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_66
timestamp 1623529830
transform 1 0 7176 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_78
timestamp 1623529830
transform 1 0 8280 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_87
timestamp 1623529830
transform 1 0 9108 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_99
timestamp 1623529830
transform 1 0 10212 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_111
timestamp 1623529830
transform 1 0 11316 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_123
timestamp 1623529830
transform 1 0 12420 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1623529830
transform 1 0 14260 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_135
timestamp 1623529830
transform 1 0 13524 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_144
timestamp 1623529830
transform 1 0 14352 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_156
timestamp 1623529830
transform 1 0 15456 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_168
timestamp 1623529830
transform 1 0 16560 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_180
timestamp 1623529830
transform 1 0 17664 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_192
timestamp 1623529830
transform 1 0 18768 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1623529830
transform 1 0 19504 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_201
timestamp 1623529830
transform 1 0 19596 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_213
timestamp 1623529830
transform 1 0 20700 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_225
timestamp 1623529830
transform 1 0 21804 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_237
timestamp 1623529830
transform 1 0 22908 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1623529830
transform 1 0 24748 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_249
timestamp 1623529830
transform 1 0 24012 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_258
timestamp 1623529830
transform 1 0 24840 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_270
timestamp 1623529830
transform 1 0 25944 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_282
timestamp 1623529830
transform 1 0 27048 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_294
timestamp 1623529830
transform 1 0 28152 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1623529830
transform 1 0 29992 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_306
timestamp 1623529830
transform 1 0 29256 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_315
timestamp 1623529830
transform 1 0 30084 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_327
timestamp 1623529830
transform 1 0 31188 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_339
timestamp 1623529830
transform 1 0 32292 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1623529830
transform 1 0 35236 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_351
timestamp 1623529830
transform 1 0 33396 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_363
timestamp 1623529830
transform 1 0 34500 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_372
timestamp 1623529830
transform 1 0 35328 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_384
timestamp 1623529830
transform 1 0 36432 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1623529830
transform -1 0 38824 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_396
timestamp 1623529830
transform 1 0 37536 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_404
timestamp 1623529830
transform 1 0 38272 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1623529830
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1623529830
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1623529830
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1623529830
transform 1 0 3588 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1623529830
transform 1 0 4692 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1623529830
transform 1 0 6348 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_51
timestamp 1623529830
transform 1 0 5796 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_58
timestamp 1623529830
transform 1 0 6440 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_70
timestamp 1623529830
transform 1 0 7544 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_82
timestamp 1623529830
transform 1 0 8648 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_94
timestamp 1623529830
transform 1 0 9752 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_106
timestamp 1623529830
transform 1 0 10856 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1623529830
transform 1 0 11592 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_115
timestamp 1623529830
transform 1 0 11684 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_127
timestamp 1623529830
transform 1 0 12788 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_139
timestamp 1623529830
transform 1 0 13892 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_151
timestamp 1623529830
transform 1 0 14996 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1623529830
transform 1 0 16836 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_163
timestamp 1623529830
transform 1 0 16100 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_172
timestamp 1623529830
transform 1 0 16928 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_184
timestamp 1623529830
transform 1 0 18032 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_196
timestamp 1623529830
transform 1 0 19136 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_208
timestamp 1623529830
transform 1 0 20240 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1623529830
transform 1 0 22080 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_220
timestamp 1623529830
transform 1 0 21344 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_229
timestamp 1623529830
transform 1 0 22172 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_241
timestamp 1623529830
transform 1 0 23276 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_253
timestamp 1623529830
transform 1 0 24380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_265
timestamp 1623529830
transform 1 0 25484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_277
timestamp 1623529830
transform 1 0 26588 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1623529830
transform 1 0 27324 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_286
timestamp 1623529830
transform 1 0 27416 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_298
timestamp 1623529830
transform 1 0 28520 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_310
timestamp 1623529830
transform 1 0 29624 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_322
timestamp 1623529830
transform 1 0 30728 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1623529830
transform 1 0 32568 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_334
timestamp 1623529830
transform 1 0 31832 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_343
timestamp 1623529830
transform 1 0 32660 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_355
timestamp 1623529830
transform 1 0 33764 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_367
timestamp 1623529830
transform 1 0 34868 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_379
timestamp 1623529830
transform 1 0 35972 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_391
timestamp 1623529830
transform 1 0 37076 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1623529830
transform -1 0 38824 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1623529830
transform 1 0 37812 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_400
timestamp 1623529830
transform 1 0 37904 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_406
timestamp 1623529830
transform 1 0 38456 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1623529830
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1623529830
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1623529830
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1623529830
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1623529830
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1623529830
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1623529830
transform 1 0 3772 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_27
timestamp 1623529830
transform 1 0 3588 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_30
timestamp 1623529830
transform 1 0 3864 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_42
timestamp 1623529830
transform 1 0 4968 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1623529830
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1623529830
transform 1 0 4692 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1623529830
transform 1 0 6348 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_54
timestamp 1623529830
transform 1 0 6072 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_51
timestamp 1623529830
transform 1 0 5796 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_58
timestamp 1623529830
transform 1 0 6440 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1623529830
transform 1 0 9016 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_66
timestamp 1623529830
transform 1 0 7176 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_78
timestamp 1623529830
transform 1 0 8280 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_87
timestamp 1623529830
transform 1 0 9108 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_70
timestamp 1623529830
transform 1 0 7544 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_82
timestamp 1623529830
transform 1 0 8648 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_99
timestamp 1623529830
transform 1 0 10212 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_94
timestamp 1623529830
transform 1 0 9752 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_106
timestamp 1623529830
transform 1 0 10856 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1623529830
transform 1 0 11592 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_111
timestamp 1623529830
transform 1 0 11316 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_123
timestamp 1623529830
transform 1 0 12420 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_115
timestamp 1623529830
transform 1 0 11684 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_127
timestamp 1623529830
transform 1 0 12788 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1623529830
transform 1 0 14260 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_135
timestamp 1623529830
transform 1 0 13524 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_144
timestamp 1623529830
transform 1 0 14352 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_139
timestamp 1623529830
transform 1 0 13892 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_151
timestamp 1623529830
transform 1 0 14996 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1623529830
transform 1 0 16836 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_156
timestamp 1623529830
transform 1 0 15456 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_168
timestamp 1623529830
transform 1 0 16560 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_163
timestamp 1623529830
transform 1 0 16100 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_172
timestamp 1623529830
transform 1 0 16928 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_180
timestamp 1623529830
transform 1 0 17664 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_192
timestamp 1623529830
transform 1 0 18768 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_184
timestamp 1623529830
transform 1 0 18032 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_196
timestamp 1623529830
transform 1 0 19136 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1623529830
transform 1 0 19504 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_201
timestamp 1623529830
transform 1 0 19596 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_213
timestamp 1623529830
transform 1 0 20700 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_208
timestamp 1623529830
transform 1 0 20240 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1623529830
transform 1 0 22080 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_225
timestamp 1623529830
transform 1 0 21804 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_237
timestamp 1623529830
transform 1 0 22908 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_220
timestamp 1623529830
transform 1 0 21344 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_229
timestamp 1623529830
transform 1 0 22172 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1623529830
transform 1 0 24748 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_249
timestamp 1623529830
transform 1 0 24012 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_258
timestamp 1623529830
transform 1 0 24840 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_241
timestamp 1623529830
transform 1 0 23276 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_253
timestamp 1623529830
transform 1 0 24380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_270
timestamp 1623529830
transform 1 0 25944 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_282
timestamp 1623529830
transform 1 0 27048 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_265
timestamp 1623529830
transform 1 0 25484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_277
timestamp 1623529830
transform 1 0 26588 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1623529830
transform 1 0 27324 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_294
timestamp 1623529830
transform 1 0 28152 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_286
timestamp 1623529830
transform 1 0 27416 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_298
timestamp 1623529830
transform 1 0 28520 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1623529830
transform 1 0 29992 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_306
timestamp 1623529830
transform 1 0 29256 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_315
timestamp 1623529830
transform 1 0 30084 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_327
timestamp 1623529830
transform 1 0 31188 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_310
timestamp 1623529830
transform 1 0 29624 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_322
timestamp 1623529830
transform 1 0 30728 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1623529830
transform 1 0 32568 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_339
timestamp 1623529830
transform 1 0 32292 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_334
timestamp 1623529830
transform 1 0 31832 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_343
timestamp 1623529830
transform 1 0 32660 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1623529830
transform 1 0 35236 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_351
timestamp 1623529830
transform 1 0 33396 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_363
timestamp 1623529830
transform 1 0 34500 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_355
timestamp 1623529830
transform 1 0 33764 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_367
timestamp 1623529830
transform 1 0 34868 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_372
timestamp 1623529830
transform 1 0 35328 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_384
timestamp 1623529830
transform 1 0 36432 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_379
timestamp 1623529830
transform 1 0 35972 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_391
timestamp 1623529830
transform 1 0 37076 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1623529830
transform -1 0 38824 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1623529830
transform -1 0 38824 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1623529830
transform 1 0 37812 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_396
timestamp 1623529830
transform 1 0 37536 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_404
timestamp 1623529830
transform 1 0 38272 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_400
timestamp 1623529830
transform 1 0 37904 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_406
timestamp 1623529830
transform 1 0 38456 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1623529830
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1623529830
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1623529830
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1623529830
transform 1 0 3772 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_27
timestamp 1623529830
transform 1 0 3588 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_30
timestamp 1623529830
transform 1 0 3864 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_42
timestamp 1623529830
transform 1 0 4968 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_54
timestamp 1623529830
transform 1 0 6072 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1623529830
transform 1 0 9016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_66
timestamp 1623529830
transform 1 0 7176 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_78
timestamp 1623529830
transform 1 0 8280 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_87
timestamp 1623529830
transform 1 0 9108 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_99
timestamp 1623529830
transform 1 0 10212 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_111
timestamp 1623529830
transform 1 0 11316 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_123
timestamp 1623529830
transform 1 0 12420 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1623529830
transform 1 0 14260 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_135
timestamp 1623529830
transform 1 0 13524 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_144
timestamp 1623529830
transform 1 0 14352 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_156
timestamp 1623529830
transform 1 0 15456 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_168
timestamp 1623529830
transform 1 0 16560 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_180
timestamp 1623529830
transform 1 0 17664 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_192
timestamp 1623529830
transform 1 0 18768 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1623529830
transform 1 0 19504 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_201
timestamp 1623529830
transform 1 0 19596 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_213
timestamp 1623529830
transform 1 0 20700 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_225
timestamp 1623529830
transform 1 0 21804 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_237
timestamp 1623529830
transform 1 0 22908 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1623529830
transform 1 0 24748 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_249
timestamp 1623529830
transform 1 0 24012 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_258
timestamp 1623529830
transform 1 0 24840 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_270
timestamp 1623529830
transform 1 0 25944 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_282
timestamp 1623529830
transform 1 0 27048 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_294
timestamp 1623529830
transform 1 0 28152 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1623529830
transform 1 0 29992 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_306
timestamp 1623529830
transform 1 0 29256 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_315
timestamp 1623529830
transform 1 0 30084 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_327
timestamp 1623529830
transform 1 0 31188 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_339
timestamp 1623529830
transform 1 0 32292 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1623529830
transform 1 0 35236 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_351
timestamp 1623529830
transform 1 0 33396 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_363
timestamp 1623529830
transform 1 0 34500 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_372
timestamp 1623529830
transform 1 0 35328 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_384
timestamp 1623529830
transform 1 0 36432 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1623529830
transform -1 0 38824 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_396
timestamp 1623529830
transform 1 0 37536 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_404
timestamp 1623529830
transform 1 0 38272 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1623529830
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1623529830
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1623529830
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1623529830
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1623529830
transform 1 0 4692 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1623529830
transform 1 0 6348 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_51
timestamp 1623529830
transform 1 0 5796 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_58
timestamp 1623529830
transform 1 0 6440 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_70
timestamp 1623529830
transform 1 0 7544 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_82
timestamp 1623529830
transform 1 0 8648 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_94
timestamp 1623529830
transform 1 0 9752 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_106
timestamp 1623529830
transform 1 0 10856 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1623529830
transform 1 0 11592 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_115
timestamp 1623529830
transform 1 0 11684 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_127
timestamp 1623529830
transform 1 0 12788 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_139
timestamp 1623529830
transform 1 0 13892 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_151
timestamp 1623529830
transform 1 0 14996 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1623529830
transform 1 0 16836 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_163
timestamp 1623529830
transform 1 0 16100 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_172
timestamp 1623529830
transform 1 0 16928 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_184
timestamp 1623529830
transform 1 0 18032 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_196
timestamp 1623529830
transform 1 0 19136 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_208
timestamp 1623529830
transform 1 0 20240 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1623529830
transform 1 0 22080 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_220
timestamp 1623529830
transform 1 0 21344 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_229
timestamp 1623529830
transform 1 0 22172 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_241
timestamp 1623529830
transform 1 0 23276 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_253
timestamp 1623529830
transform 1 0 24380 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_265
timestamp 1623529830
transform 1 0 25484 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_277
timestamp 1623529830
transform 1 0 26588 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1623529830
transform 1 0 27324 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_286
timestamp 1623529830
transform 1 0 27416 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_298
timestamp 1623529830
transform 1 0 28520 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_310
timestamp 1623529830
transform 1 0 29624 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_322
timestamp 1623529830
transform 1 0 30728 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1623529830
transform 1 0 32568 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_334
timestamp 1623529830
transform 1 0 31832 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_343
timestamp 1623529830
transform 1 0 32660 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_355
timestamp 1623529830
transform 1 0 33764 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_367
timestamp 1623529830
transform 1 0 34868 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_379
timestamp 1623529830
transform 1 0 35972 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_391
timestamp 1623529830
transform 1 0 37076 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1623529830
transform -1 0 38824 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1623529830
transform 1 0 37812 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_400
timestamp 1623529830
transform 1 0 37904 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_406
timestamp 1623529830
transform 1 0 38456 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1623529830
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1623529830
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1623529830
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1623529830
transform 1 0 3772 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_27
timestamp 1623529830
transform 1 0 3588 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_30
timestamp 1623529830
transform 1 0 3864 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_42
timestamp 1623529830
transform 1 0 4968 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_54
timestamp 1623529830
transform 1 0 6072 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1623529830
transform 1 0 9016 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_66
timestamp 1623529830
transform 1 0 7176 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_78
timestamp 1623529830
transform 1 0 8280 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_87
timestamp 1623529830
transform 1 0 9108 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_99
timestamp 1623529830
transform 1 0 10212 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_111
timestamp 1623529830
transform 1 0 11316 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_123
timestamp 1623529830
transform 1 0 12420 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1623529830
transform 1 0 14260 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_135
timestamp 1623529830
transform 1 0 13524 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_144
timestamp 1623529830
transform 1 0 14352 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_156
timestamp 1623529830
transform 1 0 15456 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_168
timestamp 1623529830
transform 1 0 16560 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_180
timestamp 1623529830
transform 1 0 17664 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_192
timestamp 1623529830
transform 1 0 18768 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1623529830
transform 1 0 19504 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_201
timestamp 1623529830
transform 1 0 19596 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_213
timestamp 1623529830
transform 1 0 20700 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_225
timestamp 1623529830
transform 1 0 21804 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_237
timestamp 1623529830
transform 1 0 22908 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1623529830
transform 1 0 24748 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_249
timestamp 1623529830
transform 1 0 24012 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_258
timestamp 1623529830
transform 1 0 24840 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_270
timestamp 1623529830
transform 1 0 25944 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_282
timestamp 1623529830
transform 1 0 27048 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_294
timestamp 1623529830
transform 1 0 28152 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1623529830
transform 1 0 29992 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_306
timestamp 1623529830
transform 1 0 29256 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_315
timestamp 1623529830
transform 1 0 30084 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_327
timestamp 1623529830
transform 1 0 31188 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_339
timestamp 1623529830
transform 1 0 32292 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1623529830
transform 1 0 35236 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_351
timestamp 1623529830
transform 1 0 33396 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_363
timestamp 1623529830
transform 1 0 34500 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_372
timestamp 1623529830
transform 1 0 35328 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_384
timestamp 1623529830
transform 1 0 36432 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1623529830
transform -1 0 38824 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_396
timestamp 1623529830
transform 1 0 37536 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_404
timestamp 1623529830
transform 1 0 38272 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1623529830
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1623529830
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1623529830
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1623529830
transform 1 0 3588 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1623529830
transform 1 0 4692 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1623529830
transform 1 0 6348 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_51
timestamp 1623529830
transform 1 0 5796 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_58
timestamp 1623529830
transform 1 0 6440 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_70
timestamp 1623529830
transform 1 0 7544 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_82
timestamp 1623529830
transform 1 0 8648 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_94
timestamp 1623529830
transform 1 0 9752 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_106
timestamp 1623529830
transform 1 0 10856 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1623529830
transform 1 0 11592 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_115
timestamp 1623529830
transform 1 0 11684 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_127
timestamp 1623529830
transform 1 0 12788 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_139
timestamp 1623529830
transform 1 0 13892 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_151
timestamp 1623529830
transform 1 0 14996 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1623529830
transform 1 0 16836 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_163
timestamp 1623529830
transform 1 0 16100 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_172
timestamp 1623529830
transform 1 0 16928 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_184
timestamp 1623529830
transform 1 0 18032 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_196
timestamp 1623529830
transform 1 0 19136 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_208
timestamp 1623529830
transform 1 0 20240 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1623529830
transform 1 0 22080 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_220
timestamp 1623529830
transform 1 0 21344 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_229
timestamp 1623529830
transform 1 0 22172 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_241
timestamp 1623529830
transform 1 0 23276 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_253
timestamp 1623529830
transform 1 0 24380 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_265
timestamp 1623529830
transform 1 0 25484 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_277
timestamp 1623529830
transform 1 0 26588 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1623529830
transform 1 0 27324 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_286
timestamp 1623529830
transform 1 0 27416 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_298
timestamp 1623529830
transform 1 0 28520 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_310
timestamp 1623529830
transform 1 0 29624 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_322
timestamp 1623529830
transform 1 0 30728 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1623529830
transform 1 0 32568 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_334
timestamp 1623529830
transform 1 0 31832 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_343
timestamp 1623529830
transform 1 0 32660 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_355
timestamp 1623529830
transform 1 0 33764 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_367
timestamp 1623529830
transform 1 0 34868 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_379
timestamp 1623529830
transform 1 0 35972 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_391
timestamp 1623529830
transform 1 0 37076 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1623529830
transform -1 0 38824 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1623529830
transform 1 0 37812 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_400
timestamp 1623529830
transform 1 0 37904 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_406
timestamp 1623529830
transform 1 0 38456 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1623529830
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1623529830
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1623529830
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1623529830
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1623529830
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1623529830
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1623529830
transform 1 0 3772 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_27
timestamp 1623529830
transform 1 0 3588 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_30
timestamp 1623529830
transform 1 0 3864 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_42
timestamp 1623529830
transform 1 0 4968 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1623529830
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1623529830
transform 1 0 4692 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1623529830
transform 1 0 6348 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_54
timestamp 1623529830
transform 1 0 6072 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_51
timestamp 1623529830
transform 1 0 5796 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_58
timestamp 1623529830
transform 1 0 6440 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1623529830
transform 1 0 9016 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_66
timestamp 1623529830
transform 1 0 7176 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_78
timestamp 1623529830
transform 1 0 8280 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_87
timestamp 1623529830
transform 1 0 9108 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_70
timestamp 1623529830
transform 1 0 7544 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_82
timestamp 1623529830
transform 1 0 8648 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_99
timestamp 1623529830
transform 1 0 10212 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_94
timestamp 1623529830
transform 1 0 9752 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_106
timestamp 1623529830
transform 1 0 10856 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1623529830
transform 1 0 11592 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_111
timestamp 1623529830
transform 1 0 11316 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_123
timestamp 1623529830
transform 1 0 12420 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_115
timestamp 1623529830
transform 1 0 11684 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_127
timestamp 1623529830
transform 1 0 12788 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1623529830
transform 1 0 14260 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_135
timestamp 1623529830
transform 1 0 13524 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_144
timestamp 1623529830
transform 1 0 14352 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_139
timestamp 1623529830
transform 1 0 13892 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_151
timestamp 1623529830
transform 1 0 14996 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1623529830
transform 1 0 16836 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_156
timestamp 1623529830
transform 1 0 15456 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_168
timestamp 1623529830
transform 1 0 16560 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_163
timestamp 1623529830
transform 1 0 16100 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_172
timestamp 1623529830
transform 1 0 16928 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_180
timestamp 1623529830
transform 1 0 17664 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_192
timestamp 1623529830
transform 1 0 18768 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_184
timestamp 1623529830
transform 1 0 18032 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_196
timestamp 1623529830
transform 1 0 19136 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1623529830
transform 1 0 19504 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_201
timestamp 1623529830
transform 1 0 19596 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_213
timestamp 1623529830
transform 1 0 20700 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_208
timestamp 1623529830
transform 1 0 20240 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1623529830
transform 1 0 22080 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_225
timestamp 1623529830
transform 1 0 21804 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_237
timestamp 1623529830
transform 1 0 22908 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_220
timestamp 1623529830
transform 1 0 21344 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_229
timestamp 1623529830
transform 1 0 22172 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1623529830
transform 1 0 24748 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_249
timestamp 1623529830
transform 1 0 24012 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_258
timestamp 1623529830
transform 1 0 24840 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_241
timestamp 1623529830
transform 1 0 23276 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_253
timestamp 1623529830
transform 1 0 24380 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_270
timestamp 1623529830
transform 1 0 25944 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_282
timestamp 1623529830
transform 1 0 27048 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_265
timestamp 1623529830
transform 1 0 25484 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_277
timestamp 1623529830
transform 1 0 26588 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1623529830
transform 1 0 27324 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_294
timestamp 1623529830
transform 1 0 28152 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_286
timestamp 1623529830
transform 1 0 27416 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_298
timestamp 1623529830
transform 1 0 28520 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1623529830
transform 1 0 29992 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_306
timestamp 1623529830
transform 1 0 29256 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_315
timestamp 1623529830
transform 1 0 30084 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_327
timestamp 1623529830
transform 1 0 31188 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_310
timestamp 1623529830
transform 1 0 29624 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_322
timestamp 1623529830
transform 1 0 30728 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1623529830
transform 1 0 32568 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_339
timestamp 1623529830
transform 1 0 32292 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_334
timestamp 1623529830
transform 1 0 31832 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_343
timestamp 1623529830
transform 1 0 32660 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1623529830
transform 1 0 35236 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_351
timestamp 1623529830
transform 1 0 33396 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_363
timestamp 1623529830
transform 1 0 34500 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_355
timestamp 1623529830
transform 1 0 33764 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_367
timestamp 1623529830
transform 1 0 34868 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_372
timestamp 1623529830
transform 1 0 35328 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_384
timestamp 1623529830
transform 1 0 36432 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_379
timestamp 1623529830
transform 1 0 35972 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_391
timestamp 1623529830
transform 1 0 37076 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1623529830
transform -1 0 38824 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1623529830
transform -1 0 38824 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1623529830
transform 1 0 37812 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_396
timestamp 1623529830
transform 1 0 37536 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_404
timestamp 1623529830
transform 1 0 38272 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_400
timestamp 1623529830
transform 1 0 37904 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_406
timestamp 1623529830
transform 1 0 38456 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1623529830
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1623529830
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1623529830
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1623529830
transform 1 0 3772 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_27
timestamp 1623529830
transform 1 0 3588 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_30
timestamp 1623529830
transform 1 0 3864 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_42
timestamp 1623529830
transform 1 0 4968 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_54
timestamp 1623529830
transform 1 0 6072 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1623529830
transform 1 0 9016 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_66
timestamp 1623529830
transform 1 0 7176 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_78
timestamp 1623529830
transform 1 0 8280 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_87
timestamp 1623529830
transform 1 0 9108 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_99
timestamp 1623529830
transform 1 0 10212 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_111
timestamp 1623529830
transform 1 0 11316 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_123
timestamp 1623529830
transform 1 0 12420 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1623529830
transform 1 0 14260 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_135
timestamp 1623529830
transform 1 0 13524 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_144
timestamp 1623529830
transform 1 0 14352 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_156
timestamp 1623529830
transform 1 0 15456 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_168
timestamp 1623529830
transform 1 0 16560 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_180
timestamp 1623529830
transform 1 0 17664 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_192
timestamp 1623529830
transform 1 0 18768 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1623529830
transform 1 0 19504 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_201
timestamp 1623529830
transform 1 0 19596 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_213
timestamp 1623529830
transform 1 0 20700 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_225
timestamp 1623529830
transform 1 0 21804 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_237
timestamp 1623529830
transform 1 0 22908 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1623529830
transform 1 0 24748 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_249
timestamp 1623529830
transform 1 0 24012 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_258
timestamp 1623529830
transform 1 0 24840 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_270
timestamp 1623529830
transform 1 0 25944 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_282
timestamp 1623529830
transform 1 0 27048 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_294
timestamp 1623529830
transform 1 0 28152 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1623529830
transform 1 0 29992 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_306
timestamp 1623529830
transform 1 0 29256 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_315
timestamp 1623529830
transform 1 0 30084 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_327
timestamp 1623529830
transform 1 0 31188 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_339
timestamp 1623529830
transform 1 0 32292 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1623529830
transform 1 0 35236 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_351
timestamp 1623529830
transform 1 0 33396 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_363
timestamp 1623529830
transform 1 0 34500 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_372
timestamp 1623529830
transform 1 0 35328 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_384
timestamp 1623529830
transform 1 0 36432 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1623529830
transform -1 0 38824 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_396
timestamp 1623529830
transform 1 0 37536 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_404
timestamp 1623529830
transform 1 0 38272 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1623529830
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1623529830
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1623529830
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1623529830
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1623529830
transform 1 0 4692 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1623529830
transform 1 0 6348 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_51
timestamp 1623529830
transform 1 0 5796 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_58
timestamp 1623529830
transform 1 0 6440 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_70
timestamp 1623529830
transform 1 0 7544 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_82
timestamp 1623529830
transform 1 0 8648 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_94
timestamp 1623529830
transform 1 0 9752 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_106
timestamp 1623529830
transform 1 0 10856 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1623529830
transform 1 0 11592 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_115
timestamp 1623529830
transform 1 0 11684 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_127
timestamp 1623529830
transform 1 0 12788 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_139
timestamp 1623529830
transform 1 0 13892 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_151
timestamp 1623529830
transform 1 0 14996 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1623529830
transform 1 0 16836 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_163
timestamp 1623529830
transform 1 0 16100 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_172
timestamp 1623529830
transform 1 0 16928 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_184
timestamp 1623529830
transform 1 0 18032 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_196
timestamp 1623529830
transform 1 0 19136 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_208
timestamp 1623529830
transform 1 0 20240 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1623529830
transform 1 0 22080 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_220
timestamp 1623529830
transform 1 0 21344 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_229
timestamp 1623529830
transform 1 0 22172 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_241
timestamp 1623529830
transform 1 0 23276 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_253
timestamp 1623529830
transform 1 0 24380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_265
timestamp 1623529830
transform 1 0 25484 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_277
timestamp 1623529830
transform 1 0 26588 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1623529830
transform 1 0 27324 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_286
timestamp 1623529830
transform 1 0 27416 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_298
timestamp 1623529830
transform 1 0 28520 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_310
timestamp 1623529830
transform 1 0 29624 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_322
timestamp 1623529830
transform 1 0 30728 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1623529830
transform 1 0 32568 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_334
timestamp 1623529830
transform 1 0 31832 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_343
timestamp 1623529830
transform 1 0 32660 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_355
timestamp 1623529830
transform 1 0 33764 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_367
timestamp 1623529830
transform 1 0 34868 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_379
timestamp 1623529830
transform 1 0 35972 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_391
timestamp 1623529830
transform 1 0 37076 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1623529830
transform -1 0 38824 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1623529830
transform 1 0 37812 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_400
timestamp 1623529830
transform 1 0 37904 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_406
timestamp 1623529830
transform 1 0 38456 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1623529830
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1623529830
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1623529830
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1623529830
transform 1 0 3772 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_27
timestamp 1623529830
transform 1 0 3588 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_30
timestamp 1623529830
transform 1 0 3864 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_42
timestamp 1623529830
transform 1 0 4968 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_54
timestamp 1623529830
transform 1 0 6072 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1623529830
transform 1 0 9016 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_66
timestamp 1623529830
transform 1 0 7176 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_78
timestamp 1623529830
transform 1 0 8280 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_87
timestamp 1623529830
transform 1 0 9108 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_99
timestamp 1623529830
transform 1 0 10212 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_111
timestamp 1623529830
transform 1 0 11316 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_123
timestamp 1623529830
transform 1 0 12420 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1623529830
transform 1 0 14260 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_135
timestamp 1623529830
transform 1 0 13524 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_144
timestamp 1623529830
transform 1 0 14352 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_156
timestamp 1623529830
transform 1 0 15456 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_168
timestamp 1623529830
transform 1 0 16560 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_180
timestamp 1623529830
transform 1 0 17664 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_192
timestamp 1623529830
transform 1 0 18768 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1623529830
transform 1 0 19504 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_201
timestamp 1623529830
transform 1 0 19596 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_213
timestamp 1623529830
transform 1 0 20700 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_225
timestamp 1623529830
transform 1 0 21804 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_237
timestamp 1623529830
transform 1 0 22908 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1623529830
transform 1 0 24748 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_249
timestamp 1623529830
transform 1 0 24012 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_258
timestamp 1623529830
transform 1 0 24840 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_270
timestamp 1623529830
transform 1 0 25944 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_282
timestamp 1623529830
transform 1 0 27048 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_294
timestamp 1623529830
transform 1 0 28152 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1623529830
transform 1 0 29992 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_306
timestamp 1623529830
transform 1 0 29256 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_315
timestamp 1623529830
transform 1 0 30084 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_327
timestamp 1623529830
transform 1 0 31188 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_339
timestamp 1623529830
transform 1 0 32292 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1623529830
transform 1 0 35236 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_351
timestamp 1623529830
transform 1 0 33396 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_363
timestamp 1623529830
transform 1 0 34500 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_372
timestamp 1623529830
transform 1 0 35328 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_384
timestamp 1623529830
transform 1 0 36432 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1623529830
transform -1 0 38824 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_396
timestamp 1623529830
transform 1 0 37536 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_404
timestamp 1623529830
transform 1 0 38272 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1623529830
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1623529830
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1623529830
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1623529830
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1623529830
transform 1 0 4692 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1623529830
transform 1 0 6348 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_51
timestamp 1623529830
transform 1 0 5796 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_58
timestamp 1623529830
transform 1 0 6440 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_70
timestamp 1623529830
transform 1 0 7544 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_82
timestamp 1623529830
transform 1 0 8648 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_94
timestamp 1623529830
transform 1 0 9752 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_106
timestamp 1623529830
transform 1 0 10856 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1623529830
transform 1 0 11592 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_115
timestamp 1623529830
transform 1 0 11684 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_127
timestamp 1623529830
transform 1 0 12788 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_139
timestamp 1623529830
transform 1 0 13892 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_151
timestamp 1623529830
transform 1 0 14996 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1623529830
transform 1 0 16836 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_163
timestamp 1623529830
transform 1 0 16100 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_172
timestamp 1623529830
transform 1 0 16928 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_184
timestamp 1623529830
transform 1 0 18032 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_196
timestamp 1623529830
transform 1 0 19136 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_208
timestamp 1623529830
transform 1 0 20240 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1623529830
transform 1 0 22080 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_220
timestamp 1623529830
transform 1 0 21344 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_229
timestamp 1623529830
transform 1 0 22172 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_241
timestamp 1623529830
transform 1 0 23276 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_253
timestamp 1623529830
transform 1 0 24380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_265
timestamp 1623529830
transform 1 0 25484 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_277
timestamp 1623529830
transform 1 0 26588 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1623529830
transform 1 0 27324 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_286
timestamp 1623529830
transform 1 0 27416 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_298
timestamp 1623529830
transform 1 0 28520 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_310
timestamp 1623529830
transform 1 0 29624 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_322
timestamp 1623529830
transform 1 0 30728 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1623529830
transform 1 0 32568 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_334
timestamp 1623529830
transform 1 0 31832 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_343
timestamp 1623529830
transform 1 0 32660 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_355
timestamp 1623529830
transform 1 0 33764 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_367
timestamp 1623529830
transform 1 0 34868 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_379
timestamp 1623529830
transform 1 0 35972 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_391
timestamp 1623529830
transform 1 0 37076 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1623529830
transform -1 0 38824 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1623529830
transform 1 0 37812 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_400
timestamp 1623529830
transform 1 0 37904 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_406
timestamp 1623529830
transform 1 0 38456 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1623529830
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1623529830
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1623529830
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1623529830
transform 1 0 3772 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_27
timestamp 1623529830
transform 1 0 3588 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_30
timestamp 1623529830
transform 1 0 3864 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_42
timestamp 1623529830
transform 1 0 4968 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_54
timestamp 1623529830
transform 1 0 6072 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1623529830
transform 1 0 9016 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_66
timestamp 1623529830
transform 1 0 7176 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_78
timestamp 1623529830
transform 1 0 8280 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_87
timestamp 1623529830
transform 1 0 9108 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_99
timestamp 1623529830
transform 1 0 10212 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_111
timestamp 1623529830
transform 1 0 11316 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_123
timestamp 1623529830
transform 1 0 12420 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1623529830
transform 1 0 14260 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_135
timestamp 1623529830
transform 1 0 13524 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_144
timestamp 1623529830
transform 1 0 14352 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_156
timestamp 1623529830
transform 1 0 15456 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_168
timestamp 1623529830
transform 1 0 16560 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_180
timestamp 1623529830
transform 1 0 17664 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_192
timestamp 1623529830
transform 1 0 18768 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1623529830
transform 1 0 19504 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_201
timestamp 1623529830
transform 1 0 19596 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_213
timestamp 1623529830
transform 1 0 20700 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_225
timestamp 1623529830
transform 1 0 21804 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_237
timestamp 1623529830
transform 1 0 22908 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1623529830
transform 1 0 24748 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_249
timestamp 1623529830
transform 1 0 24012 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_258
timestamp 1623529830
transform 1 0 24840 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_270
timestamp 1623529830
transform 1 0 25944 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_282
timestamp 1623529830
transform 1 0 27048 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_294
timestamp 1623529830
transform 1 0 28152 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1623529830
transform 1 0 29992 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_306
timestamp 1623529830
transform 1 0 29256 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_315
timestamp 1623529830
transform 1 0 30084 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_327
timestamp 1623529830
transform 1 0 31188 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_339
timestamp 1623529830
transform 1 0 32292 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1623529830
transform 1 0 35236 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_351
timestamp 1623529830
transform 1 0 33396 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_363
timestamp 1623529830
transform 1 0 34500 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_372
timestamp 1623529830
transform 1 0 35328 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_384
timestamp 1623529830
transform 1 0 36432 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1623529830
transform -1 0 38824 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_396
timestamp 1623529830
transform 1 0 37536 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_404
timestamp 1623529830
transform 1 0 38272 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1623529830
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1623529830
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1623529830
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1623529830
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1623529830
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1623529830
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1623529830
transform 1 0 3772 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1623529830
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1623529830
transform 1 0 4692 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_27
timestamp 1623529830
transform 1 0 3588 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_30
timestamp 1623529830
transform 1 0 3864 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_42
timestamp 1623529830
transform 1 0 4968 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1623529830
transform 1 0 6348 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_51
timestamp 1623529830
transform 1 0 5796 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_58
timestamp 1623529830
transform 1 0 6440 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_54
timestamp 1623529830
transform 1 0 6072 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1623529830
transform 1 0 9016 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_70
timestamp 1623529830
transform 1 0 7544 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_82
timestamp 1623529830
transform 1 0 8648 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_66
timestamp 1623529830
transform 1 0 7176 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_78
timestamp 1623529830
transform 1 0 8280 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_87
timestamp 1623529830
transform 1 0 9108 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_94
timestamp 1623529830
transform 1 0 9752 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_106
timestamp 1623529830
transform 1 0 10856 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_99
timestamp 1623529830
transform 1 0 10212 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1623529830
transform 1 0 11592 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_115
timestamp 1623529830
transform 1 0 11684 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_127
timestamp 1623529830
transform 1 0 12788 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_111
timestamp 1623529830
transform 1 0 11316 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_123
timestamp 1623529830
transform 1 0 12420 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1623529830
transform 1 0 14260 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_139
timestamp 1623529830
transform 1 0 13892 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_151
timestamp 1623529830
transform 1 0 14996 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_135
timestamp 1623529830
transform 1 0 13524 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_144
timestamp 1623529830
transform 1 0 14352 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1623529830
transform 1 0 16836 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_163
timestamp 1623529830
transform 1 0 16100 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_172
timestamp 1623529830
transform 1 0 16928 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_156
timestamp 1623529830
transform 1 0 15456 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_168
timestamp 1623529830
transform 1 0 16560 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_184
timestamp 1623529830
transform 1 0 18032 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_196
timestamp 1623529830
transform 1 0 19136 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_180
timestamp 1623529830
transform 1 0 17664 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_192
timestamp 1623529830
transform 1 0 18768 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1623529830
transform 1 0 19504 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_208
timestamp 1623529830
transform 1 0 20240 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_201
timestamp 1623529830
transform 1 0 19596 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_213
timestamp 1623529830
transform 1 0 20700 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1623529830
transform 1 0 22080 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_220
timestamp 1623529830
transform 1 0 21344 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_229
timestamp 1623529830
transform 1 0 22172 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_225
timestamp 1623529830
transform 1 0 21804 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_237
timestamp 1623529830
transform 1 0 22908 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1623529830
transform 1 0 24748 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_241
timestamp 1623529830
transform 1 0 23276 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_253
timestamp 1623529830
transform 1 0 24380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_249
timestamp 1623529830
transform 1 0 24012 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_258
timestamp 1623529830
transform 1 0 24840 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_265
timestamp 1623529830
transform 1 0 25484 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_277
timestamp 1623529830
transform 1 0 26588 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_270
timestamp 1623529830
transform 1 0 25944 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_282
timestamp 1623529830
transform 1 0 27048 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1623529830
transform 1 0 27324 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_286
timestamp 1623529830
transform 1 0 27416 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_298
timestamp 1623529830
transform 1 0 28520 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_294
timestamp 1623529830
transform 1 0 28152 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1623529830
transform 1 0 29992 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_310
timestamp 1623529830
transform 1 0 29624 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_322
timestamp 1623529830
transform 1 0 30728 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_306
timestamp 1623529830
transform 1 0 29256 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_315
timestamp 1623529830
transform 1 0 30084 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_327
timestamp 1623529830
transform 1 0 31188 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1623529830
transform 1 0 32568 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_334
timestamp 1623529830
transform 1 0 31832 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_343
timestamp 1623529830
transform 1 0 32660 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_339
timestamp 1623529830
transform 1 0 32292 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1623529830
transform 1 0 35236 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_355
timestamp 1623529830
transform 1 0 33764 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_367
timestamp 1623529830
transform 1 0 34868 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_351
timestamp 1623529830
transform 1 0 33396 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_363
timestamp 1623529830
transform 1 0 34500 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_379
timestamp 1623529830
transform 1 0 35972 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_391
timestamp 1623529830
transform 1 0 37076 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_372
timestamp 1623529830
transform 1 0 35328 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_384
timestamp 1623529830
transform 1 0 36432 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1623529830
transform -1 0 38824 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1623529830
transform -1 0 38824 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1623529830
transform 1 0 37812 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_400
timestamp 1623529830
transform 1 0 37904 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_406
timestamp 1623529830
transform 1 0 38456 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_396
timestamp 1623529830
transform 1 0 37536 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_404
timestamp 1623529830
transform 1 0 38272 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1623529830
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1623529830
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1623529830
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1623529830
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1623529830
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1623529830
transform 1 0 6348 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_51
timestamp 1623529830
transform 1 0 5796 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_58
timestamp 1623529830
transform 1 0 6440 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_70
timestamp 1623529830
transform 1 0 7544 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_82
timestamp 1623529830
transform 1 0 8648 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_94
timestamp 1623529830
transform 1 0 9752 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_106
timestamp 1623529830
transform 1 0 10856 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1623529830
transform 1 0 11592 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_115
timestamp 1623529830
transform 1 0 11684 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_127
timestamp 1623529830
transform 1 0 12788 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_139
timestamp 1623529830
transform 1 0 13892 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_151
timestamp 1623529830
transform 1 0 14996 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1623529830
transform 1 0 16836 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_163
timestamp 1623529830
transform 1 0 16100 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_172
timestamp 1623529830
transform 1 0 16928 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_184
timestamp 1623529830
transform 1 0 18032 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_196
timestamp 1623529830
transform 1 0 19136 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_208
timestamp 1623529830
transform 1 0 20240 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1623529830
transform 1 0 22080 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_220
timestamp 1623529830
transform 1 0 21344 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_229
timestamp 1623529830
transform 1 0 22172 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_241
timestamp 1623529830
transform 1 0 23276 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_253
timestamp 1623529830
transform 1 0 24380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_265
timestamp 1623529830
transform 1 0 25484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_277
timestamp 1623529830
transform 1 0 26588 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1623529830
transform 1 0 27324 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_286
timestamp 1623529830
transform 1 0 27416 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_298
timestamp 1623529830
transform 1 0 28520 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_310
timestamp 1623529830
transform 1 0 29624 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_322
timestamp 1623529830
transform 1 0 30728 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1623529830
transform 1 0 32568 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_334
timestamp 1623529830
transform 1 0 31832 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_343
timestamp 1623529830
transform 1 0 32660 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_355
timestamp 1623529830
transform 1 0 33764 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_367
timestamp 1623529830
transform 1 0 34868 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_379
timestamp 1623529830
transform 1 0 35972 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_391
timestamp 1623529830
transform 1 0 37076 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1623529830
transform -1 0 38824 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1623529830
transform 1 0 37812 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_400
timestamp 1623529830
transform 1 0 37904 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_406
timestamp 1623529830
transform 1 0 38456 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1623529830
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1623529830
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1623529830
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1623529830
transform 1 0 3772 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_27
timestamp 1623529830
transform 1 0 3588 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_30
timestamp 1623529830
transform 1 0 3864 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_42
timestamp 1623529830
transform 1 0 4968 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_54
timestamp 1623529830
transform 1 0 6072 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1623529830
transform 1 0 9016 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_66
timestamp 1623529830
transform 1 0 7176 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_78
timestamp 1623529830
transform 1 0 8280 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_87
timestamp 1623529830
transform 1 0 9108 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_99
timestamp 1623529830
transform 1 0 10212 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_111
timestamp 1623529830
transform 1 0 11316 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_123
timestamp 1623529830
transform 1 0 12420 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1623529830
transform 1 0 14260 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_135
timestamp 1623529830
transform 1 0 13524 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_144
timestamp 1623529830
transform 1 0 14352 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_156
timestamp 1623529830
transform 1 0 15456 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_168
timestamp 1623529830
transform 1 0 16560 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_180
timestamp 1623529830
transform 1 0 17664 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_192
timestamp 1623529830
transform 1 0 18768 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1623529830
transform 1 0 19504 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_201
timestamp 1623529830
transform 1 0 19596 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_213
timestamp 1623529830
transform 1 0 20700 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_225
timestamp 1623529830
transform 1 0 21804 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_237
timestamp 1623529830
transform 1 0 22908 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1623529830
transform 1 0 24748 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_249
timestamp 1623529830
transform 1 0 24012 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_258
timestamp 1623529830
transform 1 0 24840 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_270
timestamp 1623529830
transform 1 0 25944 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_282
timestamp 1623529830
transform 1 0 27048 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_294
timestamp 1623529830
transform 1 0 28152 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1623529830
transform 1 0 29992 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_306
timestamp 1623529830
transform 1 0 29256 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_315
timestamp 1623529830
transform 1 0 30084 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_327
timestamp 1623529830
transform 1 0 31188 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_339
timestamp 1623529830
transform 1 0 32292 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1623529830
transform 1 0 35236 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_351
timestamp 1623529830
transform 1 0 33396 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_363
timestamp 1623529830
transform 1 0 34500 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_372
timestamp 1623529830
transform 1 0 35328 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_384
timestamp 1623529830
transform 1 0 36432 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1623529830
transform -1 0 38824 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_396
timestamp 1623529830
transform 1 0 37536 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_404
timestamp 1623529830
transform 1 0 38272 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1623529830
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1623529830
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1623529830
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1623529830
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1623529830
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1623529830
transform 1 0 6348 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_51
timestamp 1623529830
transform 1 0 5796 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_58
timestamp 1623529830
transform 1 0 6440 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_70
timestamp 1623529830
transform 1 0 7544 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_82
timestamp 1623529830
transform 1 0 8648 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_94
timestamp 1623529830
transform 1 0 9752 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_106
timestamp 1623529830
transform 1 0 10856 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1623529830
transform 1 0 11592 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_115
timestamp 1623529830
transform 1 0 11684 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_127
timestamp 1623529830
transform 1 0 12788 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_139
timestamp 1623529830
transform 1 0 13892 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_151
timestamp 1623529830
transform 1 0 14996 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1623529830
transform 1 0 16836 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_163
timestamp 1623529830
transform 1 0 16100 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_172
timestamp 1623529830
transform 1 0 16928 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_184
timestamp 1623529830
transform 1 0 18032 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_196
timestamp 1623529830
transform 1 0 19136 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_208
timestamp 1623529830
transform 1 0 20240 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1623529830
transform 1 0 22080 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_220
timestamp 1623529830
transform 1 0 21344 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_229
timestamp 1623529830
transform 1 0 22172 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_241
timestamp 1623529830
transform 1 0 23276 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_253
timestamp 1623529830
transform 1 0 24380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_265
timestamp 1623529830
transform 1 0 25484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_277
timestamp 1623529830
transform 1 0 26588 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1623529830
transform 1 0 27324 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_286
timestamp 1623529830
transform 1 0 27416 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_298
timestamp 1623529830
transform 1 0 28520 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_310
timestamp 1623529830
transform 1 0 29624 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_322
timestamp 1623529830
transform 1 0 30728 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1623529830
transform 1 0 32568 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_334
timestamp 1623529830
transform 1 0 31832 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_343
timestamp 1623529830
transform 1 0 32660 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_355
timestamp 1623529830
transform 1 0 33764 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_367
timestamp 1623529830
transform 1 0 34868 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_379
timestamp 1623529830
transform 1 0 35972 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_391
timestamp 1623529830
transform 1 0 37076 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1623529830
transform -1 0 38824 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1623529830
transform 1 0 37812 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_400
timestamp 1623529830
transform 1 0 37904 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_406
timestamp 1623529830
transform 1 0 38456 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1623529830
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1623529830
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1623529830
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1623529830
transform 1 0 3772 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_27
timestamp 1623529830
transform 1 0 3588 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_30
timestamp 1623529830
transform 1 0 3864 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_42
timestamp 1623529830
transform 1 0 4968 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1623529830
transform 1 0 6440 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_54
timestamp 1623529830
transform 1 0 6072 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_59
timestamp 1623529830
transform 1 0 6532 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1623529830
transform 1 0 9108 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_71
timestamp 1623529830
transform 1 0 7636 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_83
timestamp 1623529830
transform 1 0 8740 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_88
timestamp 1623529830
transform 1 0 9200 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_100
timestamp 1623529830
transform 1 0 10304 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1623529830
transform 1 0 11776 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_112
timestamp 1623529830
transform 1 0 11408 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_117
timestamp 1623529830
transform 1 0 11868 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_129
timestamp 1623529830
transform 1 0 12972 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1623529830
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_141
timestamp 1623529830
transform 1 0 14076 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_146
timestamp 1623529830
transform 1 0 14536 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1623529830
transform 1 0 17112 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_158
timestamp 1623529830
transform 1 0 15640 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_170
timestamp 1623529830
transform 1 0 16744 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_175
timestamp 1623529830
transform 1 0 17204 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_187
timestamp 1623529830
transform 1 0 18308 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1623529830
transform 1 0 19780 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_199
timestamp 1623529830
transform 1 0 19412 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_204
timestamp 1623529830
transform 1 0 19872 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_216
timestamp 1623529830
transform 1 0 20976 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1623529830
transform 1 0 22448 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_228
timestamp 1623529830
transform 1 0 22080 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_233
timestamp 1623529830
transform 1 0 22540 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1623529830
transform 1 0 25116 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_245
timestamp 1623529830
transform 1 0 23644 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_257
timestamp 1623529830
transform 1 0 24748 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_262
timestamp 1623529830
transform 1 0 25208 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_274
timestamp 1623529830
transform 1 0 26312 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1623529830
transform 1 0 27784 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_286
timestamp 1623529830
transform 1 0 27416 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_291
timestamp 1623529830
transform 1 0 27876 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_303
timestamp 1623529830
transform 1 0 28980 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1623529830
transform 1 0 30452 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_315
timestamp 1623529830
transform 1 0 30084 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_320
timestamp 1623529830
transform 1 0 30544 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1623529830
transform 1 0 33120 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_332
timestamp 1623529830
transform 1 0 31648 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_344
timestamp 1623529830
transform 1 0 32752 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_349
timestamp 1623529830
transform 1 0 33212 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_361
timestamp 1623529830
transform 1 0 34316 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1623529830
transform 1 0 35788 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_373
timestamp 1623529830
transform 1 0 35420 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_378
timestamp 1623529830
transform 1 0 35880 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_390
timestamp 1623529830
transform 1 0 36984 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1623529830
transform -1 0 38824 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1623529830
transform 1 0 38456 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_402
timestamp 1623529830
transform 1 0 38088 0 -1 37536
box -38 -48 406 592
<< labels >>
rlabel metal3 s 39200 20000 40000 20120 6 ARstb
port 0 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 Clk
port 1 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 LFSR0out
port 2 nsew signal tristate
rlabel metal2 s 24950 0 25006 800 6 LFSR1in
port 3 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 LFSR1out
port 4 nsew signal tristate
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 5 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 7 nsew ground bidirectional
rlabel metal4 s 35588 2176 35908 37536 6 vccd2
port 8 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 37536 6 vccd2
port 9 nsew power bidirectional
rlabel metal4 s 20228 2176 20548 37536 6 vssd2
port 10 nsew ground bidirectional
rlabel metal4 s 36248 2176 36568 37536 6 vdda1
port 11 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 37536 6 vdda1
port 12 nsew power bidirectional
rlabel metal4 s 20888 2176 21208 37536 6 vssa1
port 13 nsew ground bidirectional
rlabel metal4 s 36908 2176 37228 37536 6 vdda2
port 14 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 37536 6 vdda2
port 15 nsew power bidirectional
rlabel metal4 s 21548 2176 21868 37536 6 vssa2
port 16 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
