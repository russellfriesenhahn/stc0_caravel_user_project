magic
tech sky130A
magscale 1 2
timestamp 1624063564
<< obsli1 >>
rect 1152 2647 243360 244439
<< obsm1 >>
rect 1152 2615 243360 244471
<< metal2 >>
rect 15284 246794 15340 247594
rect 45812 246794 45868 247594
rect 76436 246794 76492 247594
rect 106964 246794 107020 247594
rect 137588 246794 137644 247594
rect 168116 246794 168172 247594
rect 198740 246794 198796 247594
rect 229268 246794 229324 247594
<< obsm2 >>
rect 1556 246738 15228 246794
rect 15396 246738 45756 246794
rect 45924 246738 76380 246794
rect 76548 246738 106908 246794
rect 107076 246738 137532 246794
rect 137700 246738 168060 246794
rect 168228 246738 198684 246794
rect 198852 246738 229212 246794
rect 229380 246738 242666 246794
rect 1556 2616 242666 246738
<< metal3 >>
rect 0 233706 800 233826
rect 0 206178 800 206298
rect 243770 206178 244570 206298
rect 0 178650 800 178770
rect 0 151122 800 151242
rect 0 123594 800 123714
rect 243770 123594 244570 123714
rect 0 96066 800 96186
rect 0 68538 800 68658
rect 0 41010 800 41130
rect 243770 41158 244570 41278
rect 0 13630 800 13750
<< obsm3 >>
rect 800 233906 243770 244455
rect 880 233626 243770 233906
rect 800 206378 243770 233626
rect 880 206098 243690 206378
rect 800 178850 243770 206098
rect 880 178570 243770 178850
rect 800 151322 243770 178570
rect 880 151042 243770 151322
rect 800 123794 243770 151042
rect 880 123514 243690 123794
rect 800 96266 243770 123514
rect 880 95986 243770 96266
rect 800 68738 243770 95986
rect 880 68458 243770 68738
rect 800 41358 243770 68458
rect 800 41210 243690 41358
rect 880 41078 243690 41210
rect 880 40930 243770 41078
rect 800 13830 243770 40930
rect 880 13550 243770 13830
rect 800 2631 243770 13550
<< metal4 >>
rect 4256 2616 4576 244470
rect 4916 2664 5236 244422
rect 5576 2664 5896 244422
rect 6236 2664 6556 244422
rect 19616 2616 19936 244470
rect 20276 2664 20596 244422
rect 20936 2664 21256 244422
rect 21596 2664 21916 244422
rect 34976 2616 35296 244470
rect 35636 2664 35956 244422
rect 36296 2664 36616 244422
rect 36956 2664 37276 244422
rect 50336 2616 50656 244470
rect 50996 2664 51316 244422
rect 51656 2664 51976 244422
rect 52316 2664 52636 244422
rect 65696 2616 66016 244470
rect 66356 2664 66676 244422
rect 67016 2664 67336 244422
rect 67676 2664 67996 244422
rect 81056 2616 81376 244470
rect 81716 2664 82036 244422
rect 82376 2664 82696 244422
rect 83036 2664 83356 244422
rect 96416 2616 96736 244470
rect 97076 2664 97396 244422
rect 97736 2664 98056 244422
rect 98396 2664 98716 244422
rect 111776 2616 112096 244470
rect 112436 2664 112756 244422
rect 113096 2664 113416 244422
rect 113756 2664 114076 244422
rect 127136 2616 127456 244470
rect 127796 2664 128116 244422
rect 128456 2664 128776 244422
rect 129116 2664 129436 244422
rect 142496 2616 142816 244470
rect 143156 2664 143476 244422
rect 143816 2664 144136 244422
rect 144476 2664 144796 244422
rect 157856 2616 158176 244470
rect 158516 2664 158836 244422
rect 159176 2664 159496 244422
rect 159836 2664 160156 244422
rect 173216 2616 173536 244470
rect 173876 2664 174196 244422
rect 174536 2664 174856 244422
rect 175196 2664 175516 244422
rect 188576 2616 188896 244470
rect 189236 2664 189556 244422
rect 189896 2664 190216 244422
rect 190556 2664 190876 244422
rect 203936 2616 204256 244470
rect 204596 2664 204916 244422
rect 205256 2664 205576 244422
rect 205916 2664 206236 244422
rect 219296 2616 219616 244470
rect 219956 2664 220276 244422
rect 220616 2664 220936 244422
rect 221276 2664 221596 244422
rect 234656 2616 234976 244470
rect 235316 2664 235636 244422
rect 235976 2664 236296 244422
rect 236636 2664 236956 244422
<< obsm4 >>
rect 46911 12177 50256 206715
rect 50736 12177 50916 206715
rect 51396 12177 51576 206715
rect 52056 12177 52236 206715
rect 52716 12177 65616 206715
rect 66096 12177 66276 206715
rect 66756 12177 66936 206715
rect 67416 12177 67596 206715
rect 68076 12177 80976 206715
rect 81456 12177 81636 206715
rect 82116 12177 82296 206715
rect 82776 12177 82956 206715
rect 83436 12177 96336 206715
rect 96816 12177 96996 206715
rect 97476 12177 97656 206715
rect 98136 12177 98316 206715
rect 98796 12177 111696 206715
rect 112176 12177 112356 206715
rect 112836 12177 113016 206715
rect 113496 12177 113676 206715
rect 114156 12177 127056 206715
rect 127536 12177 127716 206715
rect 128196 12177 128376 206715
rect 128856 12177 129036 206715
rect 129516 12177 142416 206715
rect 142896 12177 143076 206715
rect 143556 12177 143736 206715
rect 144216 12177 144396 206715
rect 144876 12177 157776 206715
rect 158256 12177 158436 206715
rect 158916 12177 159096 206715
rect 159576 12177 159756 206715
rect 160236 12177 173136 206715
rect 173616 12177 173796 206715
rect 174276 12177 174456 206715
rect 174936 12177 175116 206715
rect 175596 12177 188496 206715
rect 188976 12177 189156 206715
rect 189636 12177 189816 206715
rect 190296 12177 190476 206715
rect 190956 12177 203856 206715
rect 204336 12177 204516 206715
rect 204996 12177 205176 206715
rect 205656 12177 205836 206715
rect 206316 12177 214017 206715
<< labels >>
rlabel metal3 s 0 41010 800 41130 6 ARstb
port 1 nsew signal input
rlabel metal3 s 0 13630 800 13750 6 ClkIngress
port 2 nsew signal input
rlabel metal3 s 243770 206178 244570 206298 6 ED[0]
port 3 nsew signal output
rlabel metal3 s 243770 123594 244570 123714 6 ED[1]
port 4 nsew signal output
rlabel metal3 s 243770 41158 244570 41278 6 ED[2]
port 5 nsew signal output
rlabel metal2 s 229268 246794 229324 247594 6 ED[3]
port 6 nsew signal output
rlabel metal2 s 168116 246794 168172 247594 6 ED[4]
port 7 nsew signal output
rlabel metal2 s 137588 246794 137644 247594 6 ED[5]
port 8 nsew signal output
rlabel metal2 s 106964 246794 107020 247594 6 ED[6]
port 9 nsew signal output
rlabel metal2 s 76436 246794 76492 247594 6 ED[7]
port 10 nsew signal output
rlabel metal2 s 198740 246794 198796 247594 6 EValid
port 11 nsew signal output
rlabel metal2 s 45812 246794 45868 247594 6 ID[0]
port 12 nsew signal input
rlabel metal2 s 15284 246794 15340 247594 6 ID[1]
port 13 nsew signal input
rlabel metal3 s 0 233706 800 233826 6 ID[2]
port 14 nsew signal input
rlabel metal3 s 0 206178 800 206298 6 ID[3]
port 15 nsew signal input
rlabel metal3 s 0 151122 800 151242 6 ID[4]
port 16 nsew signal input
rlabel metal3 s 0 123594 800 123714 6 ID[5]
port 17 nsew signal input
rlabel metal3 s 0 96066 800 96186 6 ID[6]
port 18 nsew signal input
rlabel metal3 s 0 68538 800 68658 6 ID[7]
port 19 nsew signal input
rlabel metal3 s 0 178650 800 178770 6 IValid
port 20 nsew signal input
rlabel metal4 s 219296 2616 219616 244470 6 vccd1
port 21 nsew power bidirectional
rlabel metal4 s 188576 2616 188896 244470 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 157856 2616 158176 244470 6 vccd1
port 23 nsew power bidirectional
rlabel metal4 s 127136 2616 127456 244470 6 vccd1
port 24 nsew power bidirectional
rlabel metal4 s 96416 2616 96736 244470 6 vccd1
port 25 nsew power bidirectional
rlabel metal4 s 65696 2616 66016 244470 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 34976 2616 35296 244470 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 4256 2616 4576 244470 6 vccd1
port 28 nsew power bidirectional
rlabel metal4 s 234656 2616 234976 244470 6 vssd1
port 29 nsew ground bidirectional
rlabel metal4 s 203936 2616 204256 244470 6 vssd1
port 30 nsew ground bidirectional
rlabel metal4 s 173216 2616 173536 244470 6 vssd1
port 31 nsew ground bidirectional
rlabel metal4 s 142496 2616 142816 244470 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 111776 2616 112096 244470 6 vssd1
port 33 nsew ground bidirectional
rlabel metal4 s 81056 2616 81376 244470 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 50336 2616 50656 244470 6 vssd1
port 35 nsew ground bidirectional
rlabel metal4 s 19616 2616 19936 244470 6 vssd1
port 36 nsew ground bidirectional
rlabel metal4 s 219956 2664 220276 244422 6 vccd2
port 37 nsew power bidirectional
rlabel metal4 s 189236 2664 189556 244422 6 vccd2
port 38 nsew power bidirectional
rlabel metal4 s 158516 2664 158836 244422 6 vccd2
port 39 nsew power bidirectional
rlabel metal4 s 127796 2664 128116 244422 6 vccd2
port 40 nsew power bidirectional
rlabel metal4 s 97076 2664 97396 244422 6 vccd2
port 41 nsew power bidirectional
rlabel metal4 s 66356 2664 66676 244422 6 vccd2
port 42 nsew power bidirectional
rlabel metal4 s 35636 2664 35956 244422 6 vccd2
port 43 nsew power bidirectional
rlabel metal4 s 4916 2664 5236 244422 6 vccd2
port 44 nsew power bidirectional
rlabel metal4 s 235316 2664 235636 244422 6 vssd2
port 45 nsew ground bidirectional
rlabel metal4 s 204596 2664 204916 244422 6 vssd2
port 46 nsew ground bidirectional
rlabel metal4 s 173876 2664 174196 244422 6 vssd2
port 47 nsew ground bidirectional
rlabel metal4 s 143156 2664 143476 244422 6 vssd2
port 48 nsew ground bidirectional
rlabel metal4 s 112436 2664 112756 244422 6 vssd2
port 49 nsew ground bidirectional
rlabel metal4 s 81716 2664 82036 244422 6 vssd2
port 50 nsew ground bidirectional
rlabel metal4 s 50996 2664 51316 244422 6 vssd2
port 51 nsew ground bidirectional
rlabel metal4 s 20276 2664 20596 244422 6 vssd2
port 52 nsew ground bidirectional
rlabel metal4 s 220616 2664 220936 244422 6 vdda1
port 53 nsew power bidirectional
rlabel metal4 s 189896 2664 190216 244422 6 vdda1
port 54 nsew power bidirectional
rlabel metal4 s 159176 2664 159496 244422 6 vdda1
port 55 nsew power bidirectional
rlabel metal4 s 128456 2664 128776 244422 6 vdda1
port 56 nsew power bidirectional
rlabel metal4 s 97736 2664 98056 244422 6 vdda1
port 57 nsew power bidirectional
rlabel metal4 s 67016 2664 67336 244422 6 vdda1
port 58 nsew power bidirectional
rlabel metal4 s 36296 2664 36616 244422 6 vdda1
port 59 nsew power bidirectional
rlabel metal4 s 5576 2664 5896 244422 6 vdda1
port 60 nsew power bidirectional
rlabel metal4 s 235976 2664 236296 244422 6 vssa1
port 61 nsew ground bidirectional
rlabel metal4 s 205256 2664 205576 244422 6 vssa1
port 62 nsew ground bidirectional
rlabel metal4 s 174536 2664 174856 244422 6 vssa1
port 63 nsew ground bidirectional
rlabel metal4 s 143816 2664 144136 244422 6 vssa1
port 64 nsew ground bidirectional
rlabel metal4 s 113096 2664 113416 244422 6 vssa1
port 65 nsew ground bidirectional
rlabel metal4 s 82376 2664 82696 244422 6 vssa1
port 66 nsew ground bidirectional
rlabel metal4 s 51656 2664 51976 244422 6 vssa1
port 67 nsew ground bidirectional
rlabel metal4 s 20936 2664 21256 244422 6 vssa1
port 68 nsew ground bidirectional
rlabel metal4 s 221276 2664 221596 244422 6 vdda2
port 69 nsew power bidirectional
rlabel metal4 s 190556 2664 190876 244422 6 vdda2
port 70 nsew power bidirectional
rlabel metal4 s 159836 2664 160156 244422 6 vdda2
port 71 nsew power bidirectional
rlabel metal4 s 129116 2664 129436 244422 6 vdda2
port 72 nsew power bidirectional
rlabel metal4 s 98396 2664 98716 244422 6 vdda2
port 73 nsew power bidirectional
rlabel metal4 s 67676 2664 67996 244422 6 vdda2
port 74 nsew power bidirectional
rlabel metal4 s 36956 2664 37276 244422 6 vdda2
port 75 nsew power bidirectional
rlabel metal4 s 6236 2664 6556 244422 6 vdda2
port 76 nsew power bidirectional
rlabel metal4 s 236636 2664 236956 244422 6 vssa2
port 77 nsew ground bidirectional
rlabel metal4 s 205916 2664 206236 244422 6 vssa2
port 78 nsew ground bidirectional
rlabel metal4 s 175196 2664 175516 244422 6 vssa2
port 79 nsew ground bidirectional
rlabel metal4 s 144476 2664 144796 244422 6 vssa2
port 80 nsew ground bidirectional
rlabel metal4 s 113756 2664 114076 244422 6 vssa2
port 81 nsew ground bidirectional
rlabel metal4 s 83036 2664 83356 244422 6 vssa2
port 82 nsew ground bidirectional
rlabel metal4 s 52316 2664 52636 244422 6 vssa2
port 83 nsew ground bidirectional
rlabel metal4 s 21596 2664 21916 244422 6 vssa2
port 84 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 244570 247594
string LEFview TRUE
string GDS_FILE /project/openlane/stc0_core/runs/stc0_core/results/magic/stc0_core.gds
string GDS_END 79439438
string GDS_START 1577516
<< end >>

