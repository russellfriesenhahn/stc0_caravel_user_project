magic
tech sky130A
magscale 1 2
timestamp 1624023635
<< obsli1 >>
rect 1104 2159 216723 217617
<< obsm1 >>
rect 1104 2128 216735 217648
<< metal2 >>
rect 13542 219091 13598 219891
rect 40682 219091 40738 219891
rect 67914 219091 67970 219891
rect 95146 219091 95202 219891
rect 122378 219091 122434 219891
rect 149610 219091 149666 219891
rect 176842 219091 176898 219891
rect 204074 219091 204130 219891
<< obsm2 >>
rect 1306 219035 13486 219091
rect 13654 219035 40626 219091
rect 40794 219035 67858 219091
rect 68026 219035 95090 219091
rect 95258 219035 122322 219091
rect 122490 219035 149554 219091
rect 149722 219035 176786 219091
rect 176954 219035 204018 219091
rect 204186 219035 216272 219091
rect 1306 2128 216272 219035
<< metal3 >>
rect 0 207544 800 207664
rect 0 183064 800 183184
rect 216947 183200 217747 183320
rect 0 158720 800 158840
rect 0 134240 800 134360
rect 0 109760 800 109880
rect 216947 109896 217747 110016
rect 0 85416 800 85536
rect 0 60936 800 61056
rect 0 36456 800 36576
rect 216947 36592 217747 36712
rect 0 12112 800 12232
<< obsm3 >>
rect 800 207744 216947 217633
rect 880 207464 216947 207744
rect 800 183400 216947 207464
rect 800 183264 216867 183400
rect 880 183120 216867 183264
rect 880 182984 216947 183120
rect 800 158920 216947 182984
rect 880 158640 216947 158920
rect 800 134440 216947 158640
rect 880 134160 216947 134440
rect 800 110096 216947 134160
rect 800 109960 216867 110096
rect 880 109816 216867 109960
rect 880 109680 216947 109816
rect 800 85616 216947 109680
rect 880 85336 216947 85616
rect 800 61136 216947 85336
rect 880 60856 216947 61136
rect 800 36792 216947 60856
rect 800 36656 216867 36792
rect 880 36512 216867 36656
rect 880 36376 216947 36512
rect 800 12312 216947 36376
rect 880 12032 216947 12312
rect 800 2143 216947 12032
<< metal4 >>
rect 4208 2128 4528 217648
rect 4868 2176 5188 217600
rect 5528 2176 5848 217600
rect 6188 2176 6508 217600
rect 19568 2128 19888 217648
rect 20228 2176 20548 217600
rect 20888 2176 21208 217600
rect 21548 2176 21868 217600
rect 34928 2128 35248 217648
rect 35588 2176 35908 217600
rect 36248 2176 36568 217600
rect 36908 2176 37228 217600
rect 50288 2128 50608 217648
rect 50948 2176 51268 217600
rect 51608 2176 51928 217600
rect 52268 2176 52588 217600
rect 65648 2128 65968 217648
rect 66308 2176 66628 217600
rect 66968 2176 67288 217600
rect 67628 2176 67948 217600
rect 81008 2128 81328 217648
rect 81668 2176 81988 217600
rect 82328 2176 82648 217600
rect 82988 2176 83308 217600
rect 96368 2128 96688 217648
rect 97028 2176 97348 217600
rect 97688 2176 98008 217600
rect 98348 2176 98668 217600
rect 111728 2128 112048 217648
rect 112388 2176 112708 217600
rect 113048 2176 113368 217600
rect 113708 2176 114028 217600
rect 127088 2128 127408 217648
rect 127748 2176 128068 217600
rect 128408 2176 128728 217600
rect 129068 2176 129388 217600
rect 142448 2128 142768 217648
rect 143108 2176 143428 217600
rect 143768 2176 144088 217600
rect 144428 2176 144748 217600
rect 157808 2128 158128 217648
rect 158468 2176 158788 217600
rect 159128 2176 159448 217600
rect 159788 2176 160108 217600
rect 173168 2128 173488 217648
rect 173828 2176 174148 217600
rect 174488 2176 174808 217600
rect 175148 2176 175468 217600
rect 188528 2128 188848 217648
rect 189188 2176 189508 217600
rect 189848 2176 190168 217600
rect 190508 2176 190828 217600
rect 203888 2128 204208 217648
rect 204548 2176 204868 217600
rect 205208 2176 205528 217600
rect 205868 2176 206188 217600
<< obsm4 >>
rect 33179 12275 34848 210221
rect 35328 12275 35508 210221
rect 35988 12275 36168 210221
rect 36648 12275 36828 210221
rect 37308 12275 50208 210221
rect 50688 12275 50868 210221
rect 51348 12275 51528 210221
rect 52008 12275 52188 210221
rect 52668 12275 65568 210221
rect 66048 12275 66228 210221
rect 66708 12275 66888 210221
rect 67368 12275 67548 210221
rect 68028 12275 80928 210221
rect 81408 12275 81588 210221
rect 82068 12275 82248 210221
rect 82728 12275 82908 210221
rect 83388 12275 96288 210221
rect 96768 12275 96948 210221
rect 97428 12275 97608 210221
rect 98088 12275 98268 210221
rect 98748 12275 111648 210221
rect 112128 12275 112308 210221
rect 112788 12275 112968 210221
rect 113448 12275 113628 210221
rect 114108 12275 127008 210221
rect 127488 12275 127668 210221
rect 128148 12275 128328 210221
rect 128808 12275 128988 210221
rect 129468 12275 142368 210221
rect 142848 12275 143028 210221
rect 143508 12275 143688 210221
rect 144168 12275 144348 210221
rect 144828 12275 157728 210221
rect 158208 12275 158388 210221
rect 158868 12275 159048 210221
rect 159528 12275 159708 210221
rect 160188 12275 173088 210221
rect 173568 12275 173748 210221
rect 174228 12275 174408 210221
rect 174888 12275 175068 210221
rect 175548 12275 188448 210221
rect 188928 12275 189093 210221
<< labels >>
rlabel metal3 s 0 36456 800 36576 6 ARstb
port 1 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 ClkIngress
port 2 nsew signal input
rlabel metal3 s 216947 183200 217747 183320 6 ED[0]
port 3 nsew signal output
rlabel metal3 s 216947 109896 217747 110016 6 ED[1]
port 4 nsew signal output
rlabel metal3 s 216947 36592 217747 36712 6 ED[2]
port 5 nsew signal output
rlabel metal2 s 204074 219091 204130 219891 6 ED[3]
port 6 nsew signal output
rlabel metal2 s 149610 219091 149666 219891 6 ED[4]
port 7 nsew signal output
rlabel metal2 s 122378 219091 122434 219891 6 ED[5]
port 8 nsew signal output
rlabel metal2 s 95146 219091 95202 219891 6 ED[6]
port 9 nsew signal output
rlabel metal2 s 67914 219091 67970 219891 6 ED[7]
port 10 nsew signal output
rlabel metal2 s 176842 219091 176898 219891 6 EValid
port 11 nsew signal output
rlabel metal2 s 40682 219091 40738 219891 6 ID[0]
port 12 nsew signal input
rlabel metal2 s 13542 219091 13598 219891 6 ID[1]
port 13 nsew signal input
rlabel metal3 s 0 207544 800 207664 6 ID[2]
port 14 nsew signal input
rlabel metal3 s 0 183064 800 183184 6 ID[3]
port 15 nsew signal input
rlabel metal3 s 0 134240 800 134360 6 ID[4]
port 16 nsew signal input
rlabel metal3 s 0 109760 800 109880 6 ID[5]
port 17 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 ID[6]
port 18 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 ID[7]
port 19 nsew signal input
rlabel metal3 s 0 158720 800 158840 6 IValid
port 20 nsew signal input
rlabel metal4 s 188528 2128 188848 217648 6 vccd1
port 21 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 217648 6 vccd1
port 22 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 217648 6 vccd1
port 23 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 217648 6 vccd1
port 24 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 217648 6 vccd1
port 25 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 217648 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 217648 6 vccd1
port 27 nsew power bidirectional
rlabel metal4 s 203888 2128 204208 217648 6 vssd1
port 28 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 217648 6 vssd1
port 29 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 217648 6 vssd1
port 30 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 217648 6 vssd1
port 31 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 217648 6 vssd1
port 32 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 217648 6 vssd1
port 33 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 217648 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 189188 2176 189508 217600 6 vccd2
port 35 nsew power bidirectional
rlabel metal4 s 158468 2176 158788 217600 6 vccd2
port 36 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 217600 6 vccd2
port 37 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 217600 6 vccd2
port 38 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 217600 6 vccd2
port 39 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 217600 6 vccd2
port 40 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 217600 6 vccd2
port 41 nsew power bidirectional
rlabel metal4 s 204548 2176 204868 217600 6 vssd2
port 42 nsew ground bidirectional
rlabel metal4 s 173828 2176 174148 217600 6 vssd2
port 43 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 217600 6 vssd2
port 44 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 217600 6 vssd2
port 45 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 217600 6 vssd2
port 46 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 217600 6 vssd2
port 47 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 217600 6 vssd2
port 48 nsew ground bidirectional
rlabel metal4 s 189848 2176 190168 217600 6 vdda1
port 49 nsew power bidirectional
rlabel metal4 s 159128 2176 159448 217600 6 vdda1
port 50 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 217600 6 vdda1
port 51 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 217600 6 vdda1
port 52 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 217600 6 vdda1
port 53 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 217600 6 vdda1
port 54 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 217600 6 vdda1
port 55 nsew power bidirectional
rlabel metal4 s 205208 2176 205528 217600 6 vssa1
port 56 nsew ground bidirectional
rlabel metal4 s 174488 2176 174808 217600 6 vssa1
port 57 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 217600 6 vssa1
port 58 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 217600 6 vssa1
port 59 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 217600 6 vssa1
port 60 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 217600 6 vssa1
port 61 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 217600 6 vssa1
port 62 nsew ground bidirectional
rlabel metal4 s 190508 2176 190828 217600 6 vdda2
port 63 nsew power bidirectional
rlabel metal4 s 159788 2176 160108 217600 6 vdda2
port 64 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 217600 6 vdda2
port 65 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 217600 6 vdda2
port 66 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 217600 6 vdda2
port 67 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 217600 6 vdda2
port 68 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 217600 6 vdda2
port 69 nsew power bidirectional
rlabel metal4 s 205868 2176 206188 217600 6 vssa2
port 70 nsew ground bidirectional
rlabel metal4 s 175148 2176 175468 217600 6 vssa2
port 71 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 217600 6 vssa2
port 72 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 217600 6 vssa2
port 73 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 217600 6 vssa2
port 74 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 217600 6 vssa2
port 75 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 217600 6 vssa2
port 76 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 217747 219891
string LEFview TRUE
string GDS_FILE /project/openlane/stc0_core/runs/stc0_core/results/magic/stc0_core.gds
string GDS_END 81581232
string GDS_START 1455284
<< end >>

