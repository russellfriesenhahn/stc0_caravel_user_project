VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO stc0_core
  CLASS BLOCK ;
  FOREIGN stc0_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1222.850 BY 1237.970 ;
  PIN ARstb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.050 4.000 205.650 ;
    END
  END ARstb
  PIN ClkIngress
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.150 4.000 68.750 ;
    END
  END ClkIngress
  PIN ED[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1218.850 1030.890 1222.850 1031.490 ;
    END
  END ED[0]
  PIN ED[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1218.850 617.970 1222.850 618.570 ;
    END
  END ED[1]
  PIN ED[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1218.850 205.790 1222.850 206.390 ;
    END
  END ED[2]
  PIN ED[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.340 1233.970 1146.620 1237.970 ;
    END
  END ED[3]
  PIN ED[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.580 1233.970 840.860 1237.970 ;
    END
  END ED[4]
  PIN ED[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.940 1233.970 688.220 1237.970 ;
    END
  END ED[5]
  PIN ED[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.820 1233.970 535.100 1237.970 ;
    END
  END ED[6]
  PIN ED[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.180 1233.970 382.460 1237.970 ;
    END
  END ED[7]
  PIN EValid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.700 1233.970 993.980 1237.970 ;
    END
  END EValid
  PIN ID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.060 1233.970 229.340 1237.970 ;
    END
  END ID[0]
  PIN ID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.420 1233.970 76.700 1237.970 ;
    END
  END ID[1]
  PIN ID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1168.530 4.000 1169.130 ;
    END
  END ID[2]
  PIN ID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.890 4.000 1031.490 ;
    END
  END ID[3]
  PIN ID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 755.610 4.000 756.210 ;
    END
  END ID[4]
  PIN ID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.970 4.000 618.570 ;
    END
  END ID[5]
  PIN ID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.330 4.000 480.930 ;
    END
  END ID[6]
  PIN ID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.690 4.000 343.290 ;
    END
  END ID[7]
  PIN IValid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 893.250 4.000 893.850 ;
    END
  END IValid
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1096.480 13.080 1098.080 1222.350 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 942.880 13.080 944.480 1222.350 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.280 13.080 790.880 1222.350 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.680 13.080 637.280 1222.350 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 482.080 13.080 483.680 1222.350 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.480 13.080 330.080 1222.350 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.880 13.080 176.480 1222.350 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.280 13.080 22.880 1222.350 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1173.280 13.080 1174.880 1222.350 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1019.680 13.080 1021.280 1222.350 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 866.080 13.080 867.680 1222.350 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.480 13.080 714.080 1222.350 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.880 13.080 560.480 1222.350 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.280 13.080 406.880 1222.350 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.680 13.080 253.280 1222.350 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 98.080 13.080 99.680 1222.350 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1099.780 13.320 1101.380 1222.110 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 946.180 13.320 947.780 1222.110 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 792.580 13.320 794.180 1222.110 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.980 13.320 640.580 1222.110 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.380 13.320 486.980 1222.110 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.780 13.320 333.380 1222.110 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 178.180 13.320 179.780 1222.110 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.580 13.320 26.180 1222.110 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1176.580 13.320 1178.180 1222.110 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1022.980 13.320 1024.580 1222.110 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 869.380 13.320 870.980 1222.110 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 715.780 13.320 717.380 1222.110 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 562.180 13.320 563.780 1222.110 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.580 13.320 410.180 1222.110 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.980 13.320 256.580 1222.110 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.380 13.320 102.980 1222.110 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1103.080 13.320 1104.680 1222.110 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 949.480 13.320 951.080 1222.110 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 795.880 13.320 797.480 1222.110 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 642.280 13.320 643.880 1222.110 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 488.680 13.320 490.280 1222.110 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 335.080 13.320 336.680 1222.110 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.480 13.320 183.080 1222.110 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.880 13.320 29.480 1222.110 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1179.880 13.320 1181.480 1222.110 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1026.280 13.320 1027.880 1222.110 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 872.680 13.320 874.280 1222.110 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 719.080 13.320 720.680 1222.110 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 565.480 13.320 567.080 1222.110 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.880 13.320 413.480 1222.110 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.280 13.320 259.880 1222.110 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.680 13.320 106.280 1222.110 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1106.380 13.320 1107.980 1222.110 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 952.780 13.320 954.380 1222.110 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 799.180 13.320 800.780 1222.110 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 645.580 13.320 647.180 1222.110 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 491.980 13.320 493.580 1222.110 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.380 13.320 339.980 1222.110 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.780 13.320 186.380 1222.110 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 31.180 13.320 32.780 1222.110 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1183.180 13.320 1184.780 1222.110 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1029.580 13.320 1031.180 1222.110 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 875.980 13.320 877.580 1222.110 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 722.380 13.320 723.980 1222.110 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 568.780 13.320 570.380 1222.110 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 415.180 13.320 416.780 1222.110 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.580 13.320 263.180 1222.110 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.980 13.320 109.580 1222.110 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.760 13.235 1216.800 1222.195 ;
      LAYER met1 ;
        RECT 5.760 13.075 1216.800 1222.355 ;
      LAYER met2 ;
        RECT 7.780 1233.690 76.140 1233.970 ;
        RECT 76.980 1233.690 228.780 1233.970 ;
        RECT 229.620 1233.690 381.900 1233.970 ;
        RECT 382.740 1233.690 534.540 1233.970 ;
        RECT 535.380 1233.690 687.660 1233.970 ;
        RECT 688.500 1233.690 840.300 1233.970 ;
        RECT 841.140 1233.690 993.420 1233.970 ;
        RECT 994.260 1233.690 1146.060 1233.970 ;
        RECT 1146.900 1233.690 1213.330 1233.970 ;
        RECT 7.780 13.080 1213.330 1233.690 ;
      LAYER met3 ;
        RECT 4.000 1169.530 1218.850 1222.275 ;
        RECT 4.400 1168.130 1218.850 1169.530 ;
        RECT 4.000 1031.890 1218.850 1168.130 ;
        RECT 4.400 1030.490 1218.450 1031.890 ;
        RECT 4.000 894.250 1218.850 1030.490 ;
        RECT 4.400 892.850 1218.850 894.250 ;
        RECT 4.000 756.610 1218.850 892.850 ;
        RECT 4.400 755.210 1218.850 756.610 ;
        RECT 4.000 618.970 1218.850 755.210 ;
        RECT 4.400 617.570 1218.450 618.970 ;
        RECT 4.000 481.330 1218.850 617.570 ;
        RECT 4.400 479.930 1218.850 481.330 ;
        RECT 4.000 343.690 1218.850 479.930 ;
        RECT 4.400 342.290 1218.850 343.690 ;
        RECT 4.000 206.790 1218.850 342.290 ;
        RECT 4.000 206.050 1218.450 206.790 ;
        RECT 4.400 205.390 1218.450 206.050 ;
        RECT 4.400 204.650 1218.850 205.390 ;
        RECT 4.000 69.150 1218.850 204.650 ;
        RECT 4.400 67.750 1218.850 69.150 ;
        RECT 4.000 13.155 1218.850 67.750 ;
      LAYER met4 ;
        RECT 234.555 60.885 251.280 1033.575 ;
        RECT 253.680 60.885 254.580 1033.575 ;
        RECT 256.980 60.885 257.880 1033.575 ;
        RECT 260.280 60.885 261.180 1033.575 ;
        RECT 263.580 60.885 328.080 1033.575 ;
        RECT 330.480 60.885 331.380 1033.575 ;
        RECT 333.780 60.885 334.680 1033.575 ;
        RECT 337.080 60.885 337.980 1033.575 ;
        RECT 340.380 60.885 404.880 1033.575 ;
        RECT 407.280 60.885 408.180 1033.575 ;
        RECT 410.580 60.885 411.480 1033.575 ;
        RECT 413.880 60.885 414.780 1033.575 ;
        RECT 417.180 60.885 481.680 1033.575 ;
        RECT 484.080 60.885 484.980 1033.575 ;
        RECT 487.380 60.885 488.280 1033.575 ;
        RECT 490.680 60.885 491.580 1033.575 ;
        RECT 493.980 60.885 558.480 1033.575 ;
        RECT 560.880 60.885 561.780 1033.575 ;
        RECT 564.180 60.885 565.080 1033.575 ;
        RECT 567.480 60.885 568.380 1033.575 ;
        RECT 570.780 60.885 635.280 1033.575 ;
        RECT 637.680 60.885 638.580 1033.575 ;
        RECT 640.980 60.885 641.880 1033.575 ;
        RECT 644.280 60.885 645.180 1033.575 ;
        RECT 647.580 60.885 712.080 1033.575 ;
        RECT 714.480 60.885 715.380 1033.575 ;
        RECT 717.780 60.885 718.680 1033.575 ;
        RECT 721.080 60.885 721.980 1033.575 ;
        RECT 724.380 60.885 788.880 1033.575 ;
        RECT 791.280 60.885 792.180 1033.575 ;
        RECT 794.580 60.885 795.480 1033.575 ;
        RECT 797.880 60.885 798.780 1033.575 ;
        RECT 801.180 60.885 865.680 1033.575 ;
        RECT 868.080 60.885 868.980 1033.575 ;
        RECT 871.380 60.885 872.280 1033.575 ;
        RECT 874.680 60.885 875.580 1033.575 ;
        RECT 877.980 60.885 942.480 1033.575 ;
        RECT 944.880 60.885 945.780 1033.575 ;
        RECT 948.180 60.885 949.080 1033.575 ;
        RECT 951.480 60.885 952.380 1033.575 ;
        RECT 954.780 60.885 1019.280 1033.575 ;
        RECT 1021.680 60.885 1022.580 1033.575 ;
        RECT 1024.980 60.885 1025.880 1033.575 ;
        RECT 1028.280 60.885 1029.180 1033.575 ;
        RECT 1031.580 60.885 1070.085 1033.575 ;
  END
END stc0_core
END LIBRARY

